magic
tech sky130A
magscale 1 2
timestamp 1662371348
<< obsli1 >>
rect 1104 2159 11316 11985
<< obsm1 >>
rect 14 2128 11670 12016
<< metal2 >>
rect 3238 13852 3294 14652
rect 9678 13852 9734 14652
rect 18 0 74 800
rect 5814 0 5870 800
rect 11610 0 11666 800
<< obsm2 >>
rect 20 13796 3182 13852
rect 3350 13796 9622 13852
rect 9790 13796 11664 13852
rect 20 856 11664 13796
rect 130 800 5758 856
rect 5926 800 11554 856
<< metal3 >>
rect 0 12248 800 12368
rect 11708 11568 12508 11688
rect 0 6128 800 6248
rect 11708 5448 12508 5568
<< obsm3 >>
rect 880 12168 11714 12341
rect 800 11768 11714 12168
rect 800 11488 11628 11768
rect 800 6328 11714 11488
rect 880 6048 11714 6328
rect 800 5648 11714 6048
rect 800 5368 11628 5648
rect 800 2143 11714 5368
<< metal4 >>
rect 2220 2128 2540 12016
rect 3496 2128 3816 12128
rect 4773 2128 5093 12016
rect 6049 2128 6369 12128
rect 7326 2128 7646 12016
rect 8602 2128 8922 12128
rect 9879 2128 10199 12016
rect 11155 2128 11475 12128
<< metal5 >>
rect 1056 11808 11475 12128
rect 1056 10584 11364 10904
rect 1056 9360 11475 9680
rect 1056 8136 11364 8456
rect 1056 6912 11475 7232
rect 1056 5688 11364 6008
rect 1056 4464 11475 4784
rect 1056 3240 11364 3560
<< labels >>
rlabel metal2 s 18 0 74 800 6 C
port 1 nsew signal input
rlabel metal4 s 3496 2128 3816 12128 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 6049 2128 6369 12128 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 8602 2128 8922 12128 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 11155 2128 11475 12128 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 4464 11475 4784 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 6912 11475 7232 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 9360 11475 9680 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 11808 11475 12128 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 2220 2128 2540 12016 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 4773 2128 5093 12016 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 7326 2128 7646 12016 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 9879 2128 10199 12016 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 3240 11364 3560 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 5688 11364 6008 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 8136 11364 8456 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 10584 11364 10904 6 VPWR
port 3 nsew power bidirectional
rlabel metal2 s 11610 0 11666 800 6 clk
port 4 nsew signal input
rlabel metal2 s 9678 13852 9734 14652 6 light_farm[0]
port 5 nsew signal output
rlabel metal3 s 11708 11568 12508 11688 6 light_farm[1]
port 6 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 light_farm[2]
port 7 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 light_highway[0]
port 8 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 light_highway[1]
port 9 nsew signal output
rlabel metal2 s 3238 13852 3294 14652 6 light_highway[2]
port 10 nsew signal output
rlabel metal3 s 11708 5448 12508 5568 6 rst_n
port 11 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12508 14652
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 243892
string GDS_FILE /openlane/designs/iiitb_tlc/runs/RUN_2022.09.05_09.47.48/results/signoff/iiitb_tlc.magic.gds
string GDS_START 103114
<< end >>

