magic
tech sky130A
magscale 1 2
timestamp 1662371347
<< viali >>
rect 1685 11849 1719 11883
rect 4077 11849 4111 11883
rect 9965 11849 9999 11883
rect 1869 11713 1903 11747
rect 4261 11713 4295 11747
rect 9781 11713 9815 11747
rect 10517 11713 10551 11747
rect 10701 11577 10735 11611
rect 2789 11033 2823 11067
rect 2973 11033 3007 11067
rect 2881 10761 2915 10795
rect 2697 10625 2731 10659
rect 2513 10557 2547 10591
rect 4905 10557 4939 10591
rect 5181 10557 5215 10591
rect 3433 10421 3467 10455
rect 9689 9537 9723 9571
rect 3341 9469 3375 9503
rect 3709 9401 3743 9435
rect 3801 9333 3835 9367
rect 8401 9333 8435 9367
rect 5733 9129 5767 9163
rect 5549 8925 5583 8959
rect 8953 8585 8987 8619
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 10425 8381 10459 8415
rect 10701 8381 10735 8415
rect 6561 8313 6595 8347
rect 5549 8041 5583 8075
rect 9781 8041 9815 8075
rect 10057 7905 10091 7939
rect 7021 7837 7055 7871
rect 10149 7837 10183 7871
rect 4445 7497 4479 7531
rect 7849 7429 7883 7463
rect 9597 7429 9631 7463
rect 4629 7361 4663 7395
rect 10609 5865 10643 5899
rect 10793 5661 10827 5695
rect 7849 4709 7883 4743
rect 7573 4505 7607 4539
rect 8033 4437 8067 4471
rect 7849 4097 7883 4131
rect 8033 3961 8067 3995
rect 5549 3689 5583 3723
rect 9781 3689 9815 3723
rect 9137 3621 9171 3655
rect 5733 3485 5767 3519
rect 6009 3485 6043 3519
rect 6193 3485 6227 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 1777 2601 1811 2635
rect 1593 2397 1627 2431
rect 6561 2397 6595 2431
rect 6745 2261 6779 2295
<< metal1 >>
rect 1104 11994 11475 12016
rect 1104 11942 3502 11994
rect 3554 11942 3566 11994
rect 3618 11942 3630 11994
rect 3682 11942 3694 11994
rect 3746 11942 3758 11994
rect 3810 11942 6055 11994
rect 6107 11942 6119 11994
rect 6171 11942 6183 11994
rect 6235 11942 6247 11994
rect 6299 11942 6311 11994
rect 6363 11942 8608 11994
rect 8660 11942 8672 11994
rect 8724 11942 8736 11994
rect 8788 11942 8800 11994
rect 8852 11942 8864 11994
rect 8916 11942 11161 11994
rect 11213 11942 11225 11994
rect 11277 11942 11289 11994
rect 11341 11942 11353 11994
rect 11405 11942 11417 11994
rect 11469 11942 11475 11994
rect 1104 11920 11475 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 3292 11852 4077 11880
rect 3292 11840 3298 11852
rect 4065 11849 4077 11852
rect 4111 11849 4123 11883
rect 4065 11843 4123 11849
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9732 11852 9965 11880
rect 9732 11840 9738 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8352 11716 9781 11744
rect 8352 11704 8358 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 9769 11707 9827 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10686 11608 10692 11620
rect 10647 11580 10692 11608
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 1104 11450 11316 11472
rect 1104 11398 2226 11450
rect 2278 11398 2290 11450
rect 2342 11398 2354 11450
rect 2406 11398 2418 11450
rect 2470 11398 2482 11450
rect 2534 11398 4779 11450
rect 4831 11398 4843 11450
rect 4895 11398 4907 11450
rect 4959 11398 4971 11450
rect 5023 11398 5035 11450
rect 5087 11398 7332 11450
rect 7384 11398 7396 11450
rect 7448 11398 7460 11450
rect 7512 11398 7524 11450
rect 7576 11398 7588 11450
rect 7640 11398 9885 11450
rect 9937 11398 9949 11450
rect 10001 11398 10013 11450
rect 10065 11398 10077 11450
rect 10129 11398 10141 11450
rect 10193 11398 11316 11450
rect 1104 11376 11316 11398
rect 2774 11064 2780 11076
rect 2735 11036 2780 11064
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 2961 11067 3019 11073
rect 2961 11033 2973 11067
rect 3007 11064 3019 11067
rect 5626 11064 5632 11076
rect 3007 11036 5632 11064
rect 3007 11033 3019 11036
rect 2961 11027 3019 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 1104 10906 11475 10928
rect 1104 10854 3502 10906
rect 3554 10854 3566 10906
rect 3618 10854 3630 10906
rect 3682 10854 3694 10906
rect 3746 10854 3758 10906
rect 3810 10854 6055 10906
rect 6107 10854 6119 10906
rect 6171 10854 6183 10906
rect 6235 10854 6247 10906
rect 6299 10854 6311 10906
rect 6363 10854 8608 10906
rect 8660 10854 8672 10906
rect 8724 10854 8736 10906
rect 8788 10854 8800 10906
rect 8852 10854 8864 10906
rect 8916 10854 11161 10906
rect 11213 10854 11225 10906
rect 11277 10854 11289 10906
rect 11341 10854 11353 10906
rect 11405 10854 11417 10906
rect 11469 10854 11475 10906
rect 1104 10832 11475 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 7190 10792 7196 10804
rect 2915 10764 7196 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 9306 10724 9312 10736
rect 4462 10696 9312 10724
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2774 10656 2780 10668
rect 2731 10628 2780 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 4893 10591 4951 10597
rect 2547 10560 3372 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3344 10464 3372 10560
rect 4893 10557 4905 10591
rect 4939 10588 4951 10591
rect 5169 10591 5227 10597
rect 4939 10560 5120 10588
rect 4939 10557 4951 10560
rect 4893 10551 4951 10557
rect 5092 10520 5120 10560
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 5534 10588 5540 10600
rect 5215 10560 5540 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5350 10520 5356 10532
rect 5092 10492 5356 10520
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 3421 10455 3479 10461
rect 3421 10452 3433 10455
rect 3384 10424 3433 10452
rect 3384 10412 3390 10424
rect 3421 10421 3433 10424
rect 3467 10421 3479 10455
rect 3421 10415 3479 10421
rect 1104 10362 11316 10384
rect 1104 10310 2226 10362
rect 2278 10310 2290 10362
rect 2342 10310 2354 10362
rect 2406 10310 2418 10362
rect 2470 10310 2482 10362
rect 2534 10310 4779 10362
rect 4831 10310 4843 10362
rect 4895 10310 4907 10362
rect 4959 10310 4971 10362
rect 5023 10310 5035 10362
rect 5087 10310 7332 10362
rect 7384 10310 7396 10362
rect 7448 10310 7460 10362
rect 7512 10310 7524 10362
rect 7576 10310 7588 10362
rect 7640 10310 9885 10362
rect 9937 10310 9949 10362
rect 10001 10310 10013 10362
rect 10065 10310 10077 10362
rect 10129 10310 10141 10362
rect 10193 10310 11316 10362
rect 1104 10288 11316 10310
rect 1104 9818 11475 9840
rect 1104 9766 3502 9818
rect 3554 9766 3566 9818
rect 3618 9766 3630 9818
rect 3682 9766 3694 9818
rect 3746 9766 3758 9818
rect 3810 9766 6055 9818
rect 6107 9766 6119 9818
rect 6171 9766 6183 9818
rect 6235 9766 6247 9818
rect 6299 9766 6311 9818
rect 6363 9766 8608 9818
rect 8660 9766 8672 9818
rect 8724 9766 8736 9818
rect 8788 9766 8800 9818
rect 8852 9766 8864 9818
rect 8916 9766 11161 9818
rect 11213 9766 11225 9818
rect 11277 9766 11289 9818
rect 11341 9766 11353 9818
rect 11405 9766 11417 9818
rect 11469 9766 11475 9818
rect 1104 9744 11475 9766
rect 9674 9568 9680 9580
rect 9635 9540 9680 9568
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 3326 9500 3332 9512
rect 3287 9472 3332 9500
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 3697 9435 3755 9441
rect 3697 9432 3709 9435
rect 2832 9404 3709 9432
rect 2832 9392 2838 9404
rect 3697 9401 3709 9404
rect 3743 9432 3755 9435
rect 3970 9432 3976 9444
rect 3743 9404 3976 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 3786 9364 3792 9376
rect 3747 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 8386 9364 8392 9376
rect 8347 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 1104 9274 11316 9296
rect 1104 9222 2226 9274
rect 2278 9222 2290 9274
rect 2342 9222 2354 9274
rect 2406 9222 2418 9274
rect 2470 9222 2482 9274
rect 2534 9222 4779 9274
rect 4831 9222 4843 9274
rect 4895 9222 4907 9274
rect 4959 9222 4971 9274
rect 5023 9222 5035 9274
rect 5087 9222 7332 9274
rect 7384 9222 7396 9274
rect 7448 9222 7460 9274
rect 7512 9222 7524 9274
rect 7576 9222 7588 9274
rect 7640 9222 9885 9274
rect 9937 9222 9949 9274
rect 10001 9222 10013 9274
rect 10065 9222 10077 9274
rect 10129 9222 10141 9274
rect 10193 9222 11316 9274
rect 1104 9200 11316 9222
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 8294 9160 8300 9172
rect 5767 9132 8300 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 3844 8928 5549 8956
rect 3844 8916 3850 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 1104 8730 11475 8752
rect 1104 8678 3502 8730
rect 3554 8678 3566 8730
rect 3618 8678 3630 8730
rect 3682 8678 3694 8730
rect 3746 8678 3758 8730
rect 3810 8678 6055 8730
rect 6107 8678 6119 8730
rect 6171 8678 6183 8730
rect 6235 8678 6247 8730
rect 6299 8678 6311 8730
rect 6363 8678 8608 8730
rect 8660 8678 8672 8730
rect 8724 8678 8736 8730
rect 8788 8678 8800 8730
rect 8852 8678 8864 8730
rect 8916 8678 11161 8730
rect 11213 8678 11225 8730
rect 11277 8678 11289 8730
rect 11341 8678 11353 8730
rect 11405 8678 11417 8730
rect 11469 8678 11475 8730
rect 1104 8656 11475 8678
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 5684 8588 8953 8616
rect 5684 8576 5690 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 3326 8508 3332 8560
rect 3384 8548 3390 8560
rect 3384 8520 6776 8548
rect 3384 8508 3390 8520
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 6748 8489 6776 8520
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 4028 8452 6561 8480
rect 4028 8440 4034 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7834 8480 7840 8492
rect 6779 8452 7840 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6564 8412 6592 8443
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 7650 8412 7656 8424
rect 6564 8384 7656 8412
rect 7650 8372 7656 8384
rect 7708 8412 7714 8424
rect 8202 8412 8208 8424
rect 7708 8384 8208 8412
rect 7708 8372 7714 8384
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 10410 8412 10416 8424
rect 10371 8384 10416 8412
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10686 8412 10692 8424
rect 10647 8384 10692 8412
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 6546 8344 6552 8356
rect 6507 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 1104 8186 11316 8208
rect 1104 8134 2226 8186
rect 2278 8134 2290 8186
rect 2342 8134 2354 8186
rect 2406 8134 2418 8186
rect 2470 8134 2482 8186
rect 2534 8134 4779 8186
rect 4831 8134 4843 8186
rect 4895 8134 4907 8186
rect 4959 8134 4971 8186
rect 5023 8134 5035 8186
rect 5087 8134 7332 8186
rect 7384 8134 7396 8186
rect 7448 8134 7460 8186
rect 7512 8134 7524 8186
rect 7576 8134 7588 8186
rect 7640 8134 9885 8186
rect 9937 8134 9949 8186
rect 10001 8134 10013 8186
rect 10065 8134 10077 8186
rect 10129 8134 10141 8186
rect 10193 8134 11316 8186
rect 1104 8112 11316 8134
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10410 8072 10416 8084
rect 9815 8044 10416 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 8202 7896 8208 7948
rect 8260 7936 8266 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 8260 7908 10057 7936
rect 8260 7896 8266 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 8386 7868 8392 7880
rect 7055 7840 8392 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 7834 7760 7840 7812
rect 7892 7800 7898 7812
rect 10152 7800 10180 7831
rect 7892 7772 10180 7800
rect 7892 7760 7898 7772
rect 1104 7642 11475 7664
rect 1104 7590 3502 7642
rect 3554 7590 3566 7642
rect 3618 7590 3630 7642
rect 3682 7590 3694 7642
rect 3746 7590 3758 7642
rect 3810 7590 6055 7642
rect 6107 7590 6119 7642
rect 6171 7590 6183 7642
rect 6235 7590 6247 7642
rect 6299 7590 6311 7642
rect 6363 7590 8608 7642
rect 8660 7590 8672 7642
rect 8724 7590 8736 7642
rect 8788 7590 8800 7642
rect 8852 7590 8864 7642
rect 8916 7590 11161 7642
rect 11213 7590 11225 7642
rect 11277 7590 11289 7642
rect 11341 7590 11353 7642
rect 11405 7590 11417 7642
rect 11469 7590 11475 7642
rect 1104 7568 11475 7590
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4304 7500 4445 7528
rect 4304 7488 4310 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8386 7460 8392 7472
rect 7883 7432 8392 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10686 7460 10692 7472
rect 9631 7432 10692 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7392 4675 7395
rect 9766 7392 9772 7404
rect 4663 7364 9772 7392
rect 4663 7361 4675 7364
rect 4617 7355 4675 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 1104 7098 11316 7120
rect 1104 7046 2226 7098
rect 2278 7046 2290 7098
rect 2342 7046 2354 7098
rect 2406 7046 2418 7098
rect 2470 7046 2482 7098
rect 2534 7046 4779 7098
rect 4831 7046 4843 7098
rect 4895 7046 4907 7098
rect 4959 7046 4971 7098
rect 5023 7046 5035 7098
rect 5087 7046 7332 7098
rect 7384 7046 7396 7098
rect 7448 7046 7460 7098
rect 7512 7046 7524 7098
rect 7576 7046 7588 7098
rect 7640 7046 9885 7098
rect 9937 7046 9949 7098
rect 10001 7046 10013 7098
rect 10065 7046 10077 7098
rect 10129 7046 10141 7098
rect 10193 7046 11316 7098
rect 1104 7024 11316 7046
rect 1104 6554 11475 6576
rect 1104 6502 3502 6554
rect 3554 6502 3566 6554
rect 3618 6502 3630 6554
rect 3682 6502 3694 6554
rect 3746 6502 3758 6554
rect 3810 6502 6055 6554
rect 6107 6502 6119 6554
rect 6171 6502 6183 6554
rect 6235 6502 6247 6554
rect 6299 6502 6311 6554
rect 6363 6502 8608 6554
rect 8660 6502 8672 6554
rect 8724 6502 8736 6554
rect 8788 6502 8800 6554
rect 8852 6502 8864 6554
rect 8916 6502 11161 6554
rect 11213 6502 11225 6554
rect 11277 6502 11289 6554
rect 11341 6502 11353 6554
rect 11405 6502 11417 6554
rect 11469 6502 11475 6554
rect 1104 6480 11475 6502
rect 1104 6010 11316 6032
rect 1104 5958 2226 6010
rect 2278 5958 2290 6010
rect 2342 5958 2354 6010
rect 2406 5958 2418 6010
rect 2470 5958 2482 6010
rect 2534 5958 4779 6010
rect 4831 5958 4843 6010
rect 4895 5958 4907 6010
rect 4959 5958 4971 6010
rect 5023 5958 5035 6010
rect 5087 5958 7332 6010
rect 7384 5958 7396 6010
rect 7448 5958 7460 6010
rect 7512 5958 7524 6010
rect 7576 5958 7588 6010
rect 7640 5958 9885 6010
rect 9937 5958 9949 6010
rect 10001 5958 10013 6010
rect 10065 5958 10077 6010
rect 10129 5958 10141 6010
rect 10193 5958 11316 6010
rect 1104 5936 11316 5958
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 9456 5868 10609 5896
rect 9456 5856 9462 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 10597 5859 10655 5865
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 1104 5466 11475 5488
rect 1104 5414 3502 5466
rect 3554 5414 3566 5466
rect 3618 5414 3630 5466
rect 3682 5414 3694 5466
rect 3746 5414 3758 5466
rect 3810 5414 6055 5466
rect 6107 5414 6119 5466
rect 6171 5414 6183 5466
rect 6235 5414 6247 5466
rect 6299 5414 6311 5466
rect 6363 5414 8608 5466
rect 8660 5414 8672 5466
rect 8724 5414 8736 5466
rect 8788 5414 8800 5466
rect 8852 5414 8864 5466
rect 8916 5414 11161 5466
rect 11213 5414 11225 5466
rect 11277 5414 11289 5466
rect 11341 5414 11353 5466
rect 11405 5414 11417 5466
rect 11469 5414 11475 5466
rect 1104 5392 11475 5414
rect 1104 4922 11316 4944
rect 1104 4870 2226 4922
rect 2278 4870 2290 4922
rect 2342 4870 2354 4922
rect 2406 4870 2418 4922
rect 2470 4870 2482 4922
rect 2534 4870 4779 4922
rect 4831 4870 4843 4922
rect 4895 4870 4907 4922
rect 4959 4870 4971 4922
rect 5023 4870 5035 4922
rect 5087 4870 7332 4922
rect 7384 4870 7396 4922
rect 7448 4870 7460 4922
rect 7512 4870 7524 4922
rect 7576 4870 7588 4922
rect 7640 4870 9885 4922
rect 9937 4870 9949 4922
rect 10001 4870 10013 4922
rect 10065 4870 10077 4922
rect 10129 4870 10141 4922
rect 10193 4870 11316 4922
rect 1104 4848 11316 4870
rect 7834 4740 7840 4752
rect 7795 4712 7840 4740
rect 7834 4700 7840 4712
rect 7892 4700 7898 4752
rect 7561 4539 7619 4545
rect 7561 4505 7573 4539
rect 7607 4536 7619 4539
rect 7650 4536 7656 4548
rect 7607 4508 7656 4536
rect 7607 4505 7619 4508
rect 7561 4499 7619 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 9306 4468 9312 4480
rect 8067 4440 9312 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 1104 4378 11475 4400
rect 1104 4326 3502 4378
rect 3554 4326 3566 4378
rect 3618 4326 3630 4378
rect 3682 4326 3694 4378
rect 3746 4326 3758 4378
rect 3810 4326 6055 4378
rect 6107 4326 6119 4378
rect 6171 4326 6183 4378
rect 6235 4326 6247 4378
rect 6299 4326 6311 4378
rect 6363 4326 8608 4378
rect 8660 4326 8672 4378
rect 8724 4326 8736 4378
rect 8788 4326 8800 4378
rect 8852 4326 8864 4378
rect 8916 4326 11161 4378
rect 11213 4326 11225 4378
rect 11277 4326 11289 4378
rect 11341 4326 11353 4378
rect 11405 4326 11417 4378
rect 11469 4326 11475 4378
rect 1104 4304 11475 4326
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7248 4100 7849 4128
rect 7248 4088 7254 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 10502 3992 10508 4004
rect 8067 3964 10508 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 1104 3834 11316 3856
rect 1104 3782 2226 3834
rect 2278 3782 2290 3834
rect 2342 3782 2354 3834
rect 2406 3782 2418 3834
rect 2470 3782 2482 3834
rect 2534 3782 4779 3834
rect 4831 3782 4843 3834
rect 4895 3782 4907 3834
rect 4959 3782 4971 3834
rect 5023 3782 5035 3834
rect 5087 3782 7332 3834
rect 7384 3782 7396 3834
rect 7448 3782 7460 3834
rect 7512 3782 7524 3834
rect 7576 3782 7588 3834
rect 7640 3782 9885 3834
rect 9937 3782 9949 3834
rect 10001 3782 10013 3834
rect 10065 3782 10077 3834
rect 10129 3782 10141 3834
rect 10193 3782 11316 3834
rect 1104 3760 11316 3782
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5408 3692 5549 3720
rect 5408 3680 5414 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 5537 3683 5595 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 1854 3612 1860 3664
rect 1912 3652 1918 3664
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 1912 3624 9137 3652
rect 1912 3612 1918 3624
rect 9125 3621 9137 3624
rect 9171 3621 9183 3655
rect 9125 3615 9183 3621
rect 7834 3584 7840 3596
rect 5736 3556 7840 3584
rect 5736 3525 5764 3556
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 9306 3516 9312 3528
rect 6227 3488 6914 3516
rect 9267 3488 9312 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 6012 3448 6040 3479
rect 4212 3420 6040 3448
rect 6886 3448 6914 3488
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 7650 3448 7656 3460
rect 6886 3420 7656 3448
rect 4212 3408 4218 3420
rect 7650 3408 7656 3420
rect 7708 3448 7714 3460
rect 9968 3448 9996 3479
rect 7708 3420 9996 3448
rect 7708 3408 7714 3420
rect 1104 3290 11475 3312
rect 1104 3238 3502 3290
rect 3554 3238 3566 3290
rect 3618 3238 3630 3290
rect 3682 3238 3694 3290
rect 3746 3238 3758 3290
rect 3810 3238 6055 3290
rect 6107 3238 6119 3290
rect 6171 3238 6183 3290
rect 6235 3238 6247 3290
rect 6299 3238 6311 3290
rect 6363 3238 8608 3290
rect 8660 3238 8672 3290
rect 8724 3238 8736 3290
rect 8788 3238 8800 3290
rect 8852 3238 8864 3290
rect 8916 3238 11161 3290
rect 11213 3238 11225 3290
rect 11277 3238 11289 3290
rect 11341 3238 11353 3290
rect 11405 3238 11417 3290
rect 11469 3238 11475 3290
rect 1104 3216 11475 3238
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 11606 3040 11612 3052
rect 9732 3012 11612 3040
rect 9732 3000 9738 3012
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 1104 2746 11316 2768
rect 1104 2694 2226 2746
rect 2278 2694 2290 2746
rect 2342 2694 2354 2746
rect 2406 2694 2418 2746
rect 2470 2694 2482 2746
rect 2534 2694 4779 2746
rect 4831 2694 4843 2746
rect 4895 2694 4907 2746
rect 4959 2694 4971 2746
rect 5023 2694 5035 2746
rect 5087 2694 7332 2746
rect 7384 2694 7396 2746
rect 7448 2694 7460 2746
rect 7512 2694 7524 2746
rect 7576 2694 7588 2746
rect 7640 2694 9885 2746
rect 9937 2694 9949 2746
rect 10001 2694 10013 2746
rect 10065 2694 10077 2746
rect 10129 2694 10141 2746
rect 10193 2694 11316 2746
rect 1104 2672 11316 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 4154 2632 4160 2644
rect 1811 2604 4160 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 72 2400 1593 2428
rect 72 2388 78 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 1581 2391 1639 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5868 2264 6745 2292
rect 5868 2252 5874 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 1104 2202 11475 2224
rect 1104 2150 3502 2202
rect 3554 2150 3566 2202
rect 3618 2150 3630 2202
rect 3682 2150 3694 2202
rect 3746 2150 3758 2202
rect 3810 2150 6055 2202
rect 6107 2150 6119 2202
rect 6171 2150 6183 2202
rect 6235 2150 6247 2202
rect 6299 2150 6311 2202
rect 6363 2150 8608 2202
rect 8660 2150 8672 2202
rect 8724 2150 8736 2202
rect 8788 2150 8800 2202
rect 8852 2150 8864 2202
rect 8916 2150 11161 2202
rect 11213 2150 11225 2202
rect 11277 2150 11289 2202
rect 11341 2150 11353 2202
rect 11405 2150 11417 2202
rect 11469 2150 11475 2202
rect 1104 2128 11475 2150
<< via1 >>
rect 3502 11942 3554 11994
rect 3566 11942 3618 11994
rect 3630 11942 3682 11994
rect 3694 11942 3746 11994
rect 3758 11942 3810 11994
rect 6055 11942 6107 11994
rect 6119 11942 6171 11994
rect 6183 11942 6235 11994
rect 6247 11942 6299 11994
rect 6311 11942 6363 11994
rect 8608 11942 8660 11994
rect 8672 11942 8724 11994
rect 8736 11942 8788 11994
rect 8800 11942 8852 11994
rect 8864 11942 8916 11994
rect 11161 11942 11213 11994
rect 11225 11942 11277 11994
rect 11289 11942 11341 11994
rect 11353 11942 11405 11994
rect 11417 11942 11469 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 3240 11840 3292 11892
rect 9680 11840 9732 11892
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 8300 11704 8352 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10692 11611 10744 11620
rect 10692 11577 10701 11611
rect 10701 11577 10735 11611
rect 10735 11577 10744 11611
rect 10692 11568 10744 11577
rect 2226 11398 2278 11450
rect 2290 11398 2342 11450
rect 2354 11398 2406 11450
rect 2418 11398 2470 11450
rect 2482 11398 2534 11450
rect 4779 11398 4831 11450
rect 4843 11398 4895 11450
rect 4907 11398 4959 11450
rect 4971 11398 5023 11450
rect 5035 11398 5087 11450
rect 7332 11398 7384 11450
rect 7396 11398 7448 11450
rect 7460 11398 7512 11450
rect 7524 11398 7576 11450
rect 7588 11398 7640 11450
rect 9885 11398 9937 11450
rect 9949 11398 10001 11450
rect 10013 11398 10065 11450
rect 10077 11398 10129 11450
rect 10141 11398 10193 11450
rect 2780 11067 2832 11076
rect 2780 11033 2789 11067
rect 2789 11033 2823 11067
rect 2823 11033 2832 11067
rect 2780 11024 2832 11033
rect 5632 11024 5684 11076
rect 3502 10854 3554 10906
rect 3566 10854 3618 10906
rect 3630 10854 3682 10906
rect 3694 10854 3746 10906
rect 3758 10854 3810 10906
rect 6055 10854 6107 10906
rect 6119 10854 6171 10906
rect 6183 10854 6235 10906
rect 6247 10854 6299 10906
rect 6311 10854 6363 10906
rect 8608 10854 8660 10906
rect 8672 10854 8724 10906
rect 8736 10854 8788 10906
rect 8800 10854 8852 10906
rect 8864 10854 8916 10906
rect 11161 10854 11213 10906
rect 11225 10854 11277 10906
rect 11289 10854 11341 10906
rect 11353 10854 11405 10906
rect 11417 10854 11469 10906
rect 7196 10752 7248 10804
rect 9312 10684 9364 10736
rect 2780 10616 2832 10668
rect 5540 10548 5592 10600
rect 5356 10480 5408 10532
rect 3332 10412 3384 10464
rect 2226 10310 2278 10362
rect 2290 10310 2342 10362
rect 2354 10310 2406 10362
rect 2418 10310 2470 10362
rect 2482 10310 2534 10362
rect 4779 10310 4831 10362
rect 4843 10310 4895 10362
rect 4907 10310 4959 10362
rect 4971 10310 5023 10362
rect 5035 10310 5087 10362
rect 7332 10310 7384 10362
rect 7396 10310 7448 10362
rect 7460 10310 7512 10362
rect 7524 10310 7576 10362
rect 7588 10310 7640 10362
rect 9885 10310 9937 10362
rect 9949 10310 10001 10362
rect 10013 10310 10065 10362
rect 10077 10310 10129 10362
rect 10141 10310 10193 10362
rect 3502 9766 3554 9818
rect 3566 9766 3618 9818
rect 3630 9766 3682 9818
rect 3694 9766 3746 9818
rect 3758 9766 3810 9818
rect 6055 9766 6107 9818
rect 6119 9766 6171 9818
rect 6183 9766 6235 9818
rect 6247 9766 6299 9818
rect 6311 9766 6363 9818
rect 8608 9766 8660 9818
rect 8672 9766 8724 9818
rect 8736 9766 8788 9818
rect 8800 9766 8852 9818
rect 8864 9766 8916 9818
rect 11161 9766 11213 9818
rect 11225 9766 11277 9818
rect 11289 9766 11341 9818
rect 11353 9766 11405 9818
rect 11417 9766 11469 9818
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 2780 9392 2832 9444
rect 3976 9392 4028 9444
rect 3792 9367 3844 9376
rect 3792 9333 3801 9367
rect 3801 9333 3835 9367
rect 3835 9333 3844 9367
rect 3792 9324 3844 9333
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 2226 9222 2278 9274
rect 2290 9222 2342 9274
rect 2354 9222 2406 9274
rect 2418 9222 2470 9274
rect 2482 9222 2534 9274
rect 4779 9222 4831 9274
rect 4843 9222 4895 9274
rect 4907 9222 4959 9274
rect 4971 9222 5023 9274
rect 5035 9222 5087 9274
rect 7332 9222 7384 9274
rect 7396 9222 7448 9274
rect 7460 9222 7512 9274
rect 7524 9222 7576 9274
rect 7588 9222 7640 9274
rect 9885 9222 9937 9274
rect 9949 9222 10001 9274
rect 10013 9222 10065 9274
rect 10077 9222 10129 9274
rect 10141 9222 10193 9274
rect 8300 9120 8352 9172
rect 3792 8916 3844 8968
rect 3502 8678 3554 8730
rect 3566 8678 3618 8730
rect 3630 8678 3682 8730
rect 3694 8678 3746 8730
rect 3758 8678 3810 8730
rect 6055 8678 6107 8730
rect 6119 8678 6171 8730
rect 6183 8678 6235 8730
rect 6247 8678 6299 8730
rect 6311 8678 6363 8730
rect 8608 8678 8660 8730
rect 8672 8678 8724 8730
rect 8736 8678 8788 8730
rect 8800 8678 8852 8730
rect 8864 8678 8916 8730
rect 11161 8678 11213 8730
rect 11225 8678 11277 8730
rect 11289 8678 11341 8730
rect 11353 8678 11405 8730
rect 11417 8678 11469 8730
rect 5632 8576 5684 8628
rect 3332 8508 3384 8560
rect 3976 8440 4028 8492
rect 7840 8440 7892 8492
rect 9312 8440 9364 8492
rect 7656 8372 7708 8424
rect 8208 8372 8260 8424
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 2226 8134 2278 8186
rect 2290 8134 2342 8186
rect 2354 8134 2406 8186
rect 2418 8134 2470 8186
rect 2482 8134 2534 8186
rect 4779 8134 4831 8186
rect 4843 8134 4895 8186
rect 4907 8134 4959 8186
rect 4971 8134 5023 8186
rect 5035 8134 5087 8186
rect 7332 8134 7384 8186
rect 7396 8134 7448 8186
rect 7460 8134 7512 8186
rect 7524 8134 7576 8186
rect 7588 8134 7640 8186
rect 9885 8134 9937 8186
rect 9949 8134 10001 8186
rect 10013 8134 10065 8186
rect 10077 8134 10129 8186
rect 10141 8134 10193 8186
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 10416 8032 10468 8084
rect 8208 7896 8260 7948
rect 8392 7828 8444 7880
rect 7840 7760 7892 7812
rect 3502 7590 3554 7642
rect 3566 7590 3618 7642
rect 3630 7590 3682 7642
rect 3694 7590 3746 7642
rect 3758 7590 3810 7642
rect 6055 7590 6107 7642
rect 6119 7590 6171 7642
rect 6183 7590 6235 7642
rect 6247 7590 6299 7642
rect 6311 7590 6363 7642
rect 8608 7590 8660 7642
rect 8672 7590 8724 7642
rect 8736 7590 8788 7642
rect 8800 7590 8852 7642
rect 8864 7590 8916 7642
rect 11161 7590 11213 7642
rect 11225 7590 11277 7642
rect 11289 7590 11341 7642
rect 11353 7590 11405 7642
rect 11417 7590 11469 7642
rect 4252 7488 4304 7540
rect 8392 7420 8444 7472
rect 10692 7420 10744 7472
rect 9772 7352 9824 7404
rect 2226 7046 2278 7098
rect 2290 7046 2342 7098
rect 2354 7046 2406 7098
rect 2418 7046 2470 7098
rect 2482 7046 2534 7098
rect 4779 7046 4831 7098
rect 4843 7046 4895 7098
rect 4907 7046 4959 7098
rect 4971 7046 5023 7098
rect 5035 7046 5087 7098
rect 7332 7046 7384 7098
rect 7396 7046 7448 7098
rect 7460 7046 7512 7098
rect 7524 7046 7576 7098
rect 7588 7046 7640 7098
rect 9885 7046 9937 7098
rect 9949 7046 10001 7098
rect 10013 7046 10065 7098
rect 10077 7046 10129 7098
rect 10141 7046 10193 7098
rect 3502 6502 3554 6554
rect 3566 6502 3618 6554
rect 3630 6502 3682 6554
rect 3694 6502 3746 6554
rect 3758 6502 3810 6554
rect 6055 6502 6107 6554
rect 6119 6502 6171 6554
rect 6183 6502 6235 6554
rect 6247 6502 6299 6554
rect 6311 6502 6363 6554
rect 8608 6502 8660 6554
rect 8672 6502 8724 6554
rect 8736 6502 8788 6554
rect 8800 6502 8852 6554
rect 8864 6502 8916 6554
rect 11161 6502 11213 6554
rect 11225 6502 11277 6554
rect 11289 6502 11341 6554
rect 11353 6502 11405 6554
rect 11417 6502 11469 6554
rect 2226 5958 2278 6010
rect 2290 5958 2342 6010
rect 2354 5958 2406 6010
rect 2418 5958 2470 6010
rect 2482 5958 2534 6010
rect 4779 5958 4831 6010
rect 4843 5958 4895 6010
rect 4907 5958 4959 6010
rect 4971 5958 5023 6010
rect 5035 5958 5087 6010
rect 7332 5958 7384 6010
rect 7396 5958 7448 6010
rect 7460 5958 7512 6010
rect 7524 5958 7576 6010
rect 7588 5958 7640 6010
rect 9885 5958 9937 6010
rect 9949 5958 10001 6010
rect 10013 5958 10065 6010
rect 10077 5958 10129 6010
rect 10141 5958 10193 6010
rect 9404 5856 9456 5908
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 3502 5414 3554 5466
rect 3566 5414 3618 5466
rect 3630 5414 3682 5466
rect 3694 5414 3746 5466
rect 3758 5414 3810 5466
rect 6055 5414 6107 5466
rect 6119 5414 6171 5466
rect 6183 5414 6235 5466
rect 6247 5414 6299 5466
rect 6311 5414 6363 5466
rect 8608 5414 8660 5466
rect 8672 5414 8724 5466
rect 8736 5414 8788 5466
rect 8800 5414 8852 5466
rect 8864 5414 8916 5466
rect 11161 5414 11213 5466
rect 11225 5414 11277 5466
rect 11289 5414 11341 5466
rect 11353 5414 11405 5466
rect 11417 5414 11469 5466
rect 2226 4870 2278 4922
rect 2290 4870 2342 4922
rect 2354 4870 2406 4922
rect 2418 4870 2470 4922
rect 2482 4870 2534 4922
rect 4779 4870 4831 4922
rect 4843 4870 4895 4922
rect 4907 4870 4959 4922
rect 4971 4870 5023 4922
rect 5035 4870 5087 4922
rect 7332 4870 7384 4922
rect 7396 4870 7448 4922
rect 7460 4870 7512 4922
rect 7524 4870 7576 4922
rect 7588 4870 7640 4922
rect 9885 4870 9937 4922
rect 9949 4870 10001 4922
rect 10013 4870 10065 4922
rect 10077 4870 10129 4922
rect 10141 4870 10193 4922
rect 7840 4743 7892 4752
rect 7840 4709 7849 4743
rect 7849 4709 7883 4743
rect 7883 4709 7892 4743
rect 7840 4700 7892 4709
rect 7656 4496 7708 4548
rect 9312 4428 9364 4480
rect 3502 4326 3554 4378
rect 3566 4326 3618 4378
rect 3630 4326 3682 4378
rect 3694 4326 3746 4378
rect 3758 4326 3810 4378
rect 6055 4326 6107 4378
rect 6119 4326 6171 4378
rect 6183 4326 6235 4378
rect 6247 4326 6299 4378
rect 6311 4326 6363 4378
rect 8608 4326 8660 4378
rect 8672 4326 8724 4378
rect 8736 4326 8788 4378
rect 8800 4326 8852 4378
rect 8864 4326 8916 4378
rect 11161 4326 11213 4378
rect 11225 4326 11277 4378
rect 11289 4326 11341 4378
rect 11353 4326 11405 4378
rect 11417 4326 11469 4378
rect 7196 4088 7248 4140
rect 10508 3952 10560 4004
rect 2226 3782 2278 3834
rect 2290 3782 2342 3834
rect 2354 3782 2406 3834
rect 2418 3782 2470 3834
rect 2482 3782 2534 3834
rect 4779 3782 4831 3834
rect 4843 3782 4895 3834
rect 4907 3782 4959 3834
rect 4971 3782 5023 3834
rect 5035 3782 5087 3834
rect 7332 3782 7384 3834
rect 7396 3782 7448 3834
rect 7460 3782 7512 3834
rect 7524 3782 7576 3834
rect 7588 3782 7640 3834
rect 9885 3782 9937 3834
rect 9949 3782 10001 3834
rect 10013 3782 10065 3834
rect 10077 3782 10129 3834
rect 10141 3782 10193 3834
rect 5356 3680 5408 3732
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 1860 3612 1912 3664
rect 7840 3544 7892 3596
rect 9312 3519 9364 3528
rect 4160 3408 4212 3460
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 7656 3408 7708 3460
rect 3502 3238 3554 3290
rect 3566 3238 3618 3290
rect 3630 3238 3682 3290
rect 3694 3238 3746 3290
rect 3758 3238 3810 3290
rect 6055 3238 6107 3290
rect 6119 3238 6171 3290
rect 6183 3238 6235 3290
rect 6247 3238 6299 3290
rect 6311 3238 6363 3290
rect 8608 3238 8660 3290
rect 8672 3238 8724 3290
rect 8736 3238 8788 3290
rect 8800 3238 8852 3290
rect 8864 3238 8916 3290
rect 11161 3238 11213 3290
rect 11225 3238 11277 3290
rect 11289 3238 11341 3290
rect 11353 3238 11405 3290
rect 11417 3238 11469 3290
rect 9680 3000 9732 3052
rect 11612 3000 11664 3052
rect 2226 2694 2278 2746
rect 2290 2694 2342 2746
rect 2354 2694 2406 2746
rect 2418 2694 2470 2746
rect 2482 2694 2534 2746
rect 4779 2694 4831 2746
rect 4843 2694 4895 2746
rect 4907 2694 4959 2746
rect 4971 2694 5023 2746
rect 5035 2694 5087 2746
rect 7332 2694 7384 2746
rect 7396 2694 7448 2746
rect 7460 2694 7512 2746
rect 7524 2694 7576 2746
rect 7588 2694 7640 2746
rect 9885 2694 9937 2746
rect 9949 2694 10001 2746
rect 10013 2694 10065 2746
rect 10077 2694 10129 2746
rect 10141 2694 10193 2746
rect 4160 2592 4212 2644
rect 20 2388 72 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 5816 2252 5868 2304
rect 3502 2150 3554 2202
rect 3566 2150 3618 2202
rect 3630 2150 3682 2202
rect 3694 2150 3746 2202
rect 3758 2150 3810 2202
rect 6055 2150 6107 2202
rect 6119 2150 6171 2202
rect 6183 2150 6235 2202
rect 6247 2150 6299 2202
rect 6311 2150 6363 2202
rect 8608 2150 8660 2202
rect 8672 2150 8724 2202
rect 8736 2150 8788 2202
rect 8800 2150 8852 2202
rect 8864 2150 8916 2202
rect 11161 2150 11213 2202
rect 11225 2150 11277 2202
rect 11289 2150 11341 2202
rect 11353 2150 11405 2202
rect 11417 2150 11469 2202
<< metal2 >>
rect 3238 13852 3294 14652
rect 9678 13852 9734 14652
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1688 11898 1716 12271
rect 3252 11898 3280 13852
rect 3502 11996 3810 12005
rect 3502 11994 3508 11996
rect 3564 11994 3588 11996
rect 3644 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3810 11996
rect 3564 11942 3566 11994
rect 3746 11942 3748 11994
rect 3502 11940 3508 11942
rect 3564 11940 3588 11942
rect 3644 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3810 11942
rect 3502 11931 3810 11940
rect 6055 11996 6363 12005
rect 6055 11994 6061 11996
rect 6117 11994 6141 11996
rect 6197 11994 6221 11996
rect 6277 11994 6301 11996
rect 6357 11994 6363 11996
rect 6117 11942 6119 11994
rect 6299 11942 6301 11994
rect 6055 11940 6061 11942
rect 6117 11940 6141 11942
rect 6197 11940 6221 11942
rect 6277 11940 6301 11942
rect 6357 11940 6363 11942
rect 6055 11931 6363 11940
rect 8608 11996 8916 12005
rect 8608 11994 8614 11996
rect 8670 11994 8694 11996
rect 8750 11994 8774 11996
rect 8830 11994 8854 11996
rect 8910 11994 8916 11996
rect 8670 11942 8672 11994
rect 8852 11942 8854 11994
rect 8608 11940 8614 11942
rect 8670 11940 8694 11942
rect 8750 11940 8774 11942
rect 8830 11940 8854 11942
rect 8910 11940 8916 11942
rect 8608 11931 8916 11940
rect 9692 11898 9720 13852
rect 11161 11996 11469 12005
rect 11161 11994 11167 11996
rect 11223 11994 11247 11996
rect 11303 11994 11327 11996
rect 11383 11994 11407 11996
rect 11463 11994 11469 11996
rect 11223 11942 11225 11994
rect 11405 11942 11407 11994
rect 11161 11940 11167 11942
rect 11223 11940 11247 11942
rect 11303 11940 11327 11942
rect 11383 11940 11407 11942
rect 11463 11940 11469 11942
rect 11161 11931 11469 11940
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 1872 3670 1900 11698
rect 2226 11452 2534 11461
rect 2226 11450 2232 11452
rect 2288 11450 2312 11452
rect 2368 11450 2392 11452
rect 2448 11450 2472 11452
rect 2528 11450 2534 11452
rect 2288 11398 2290 11450
rect 2470 11398 2472 11450
rect 2226 11396 2232 11398
rect 2288 11396 2312 11398
rect 2368 11396 2392 11398
rect 2448 11396 2472 11398
rect 2528 11396 2534 11398
rect 2226 11387 2534 11396
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10674 2820 11018
rect 3502 10908 3810 10917
rect 3502 10906 3508 10908
rect 3564 10906 3588 10908
rect 3644 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3810 10908
rect 3564 10854 3566 10906
rect 3746 10854 3748 10906
rect 3502 10852 3508 10854
rect 3564 10852 3588 10854
rect 3644 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3810 10854
rect 3502 10843 3810 10852
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2226 10364 2534 10373
rect 2226 10362 2232 10364
rect 2288 10362 2312 10364
rect 2368 10362 2392 10364
rect 2448 10362 2472 10364
rect 2528 10362 2534 10364
rect 2288 10310 2290 10362
rect 2470 10310 2472 10362
rect 2226 10308 2232 10310
rect 2288 10308 2312 10310
rect 2368 10308 2392 10310
rect 2448 10308 2472 10310
rect 2528 10308 2534 10310
rect 2226 10299 2534 10308
rect 2792 9450 2820 10610
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 9518 3372 10406
rect 3502 9820 3810 9829
rect 3502 9818 3508 9820
rect 3564 9818 3588 9820
rect 3644 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3810 9820
rect 3564 9766 3566 9818
rect 3746 9766 3748 9818
rect 3502 9764 3508 9766
rect 3564 9764 3588 9766
rect 3644 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3810 9766
rect 3502 9755 3810 9764
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2226 9276 2534 9285
rect 2226 9274 2232 9276
rect 2288 9274 2312 9276
rect 2368 9274 2392 9276
rect 2448 9274 2472 9276
rect 2528 9274 2534 9276
rect 2288 9222 2290 9274
rect 2470 9222 2472 9274
rect 2226 9220 2232 9222
rect 2288 9220 2312 9222
rect 2368 9220 2392 9222
rect 2448 9220 2472 9222
rect 2528 9220 2534 9222
rect 2226 9211 2534 9220
rect 3344 8566 3372 9454
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 8974 3832 9318
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3502 8732 3810 8741
rect 3502 8730 3508 8732
rect 3564 8730 3588 8732
rect 3644 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3810 8732
rect 3564 8678 3566 8730
rect 3746 8678 3748 8730
rect 3502 8676 3508 8678
rect 3564 8676 3588 8678
rect 3644 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3810 8678
rect 3502 8667 3810 8676
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3988 8498 4016 9386
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 2226 8188 2534 8197
rect 2226 8186 2232 8188
rect 2288 8186 2312 8188
rect 2368 8186 2392 8188
rect 2448 8186 2472 8188
rect 2528 8186 2534 8188
rect 2288 8134 2290 8186
rect 2470 8134 2472 8186
rect 2226 8132 2232 8134
rect 2288 8132 2312 8134
rect 2368 8132 2392 8134
rect 2448 8132 2472 8134
rect 2528 8132 2534 8134
rect 2226 8123 2534 8132
rect 3502 7644 3810 7653
rect 3502 7642 3508 7644
rect 3564 7642 3588 7644
rect 3644 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3810 7644
rect 3564 7590 3566 7642
rect 3746 7590 3748 7642
rect 3502 7588 3508 7590
rect 3564 7588 3588 7590
rect 3644 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3810 7590
rect 3502 7579 3810 7588
rect 4264 7546 4292 11698
rect 4779 11452 5087 11461
rect 4779 11450 4785 11452
rect 4841 11450 4865 11452
rect 4921 11450 4945 11452
rect 5001 11450 5025 11452
rect 5081 11450 5087 11452
rect 4841 11398 4843 11450
rect 5023 11398 5025 11450
rect 4779 11396 4785 11398
rect 4841 11396 4865 11398
rect 4921 11396 4945 11398
rect 5001 11396 5025 11398
rect 5081 11396 5087 11398
rect 4779 11387 5087 11396
rect 7332 11452 7640 11461
rect 7332 11450 7338 11452
rect 7394 11450 7418 11452
rect 7474 11450 7498 11452
rect 7554 11450 7578 11452
rect 7634 11450 7640 11452
rect 7394 11398 7396 11450
rect 7576 11398 7578 11450
rect 7332 11396 7338 11398
rect 7394 11396 7418 11398
rect 7474 11396 7498 11398
rect 7554 11396 7578 11398
rect 7634 11396 7640 11398
rect 7332 11387 7640 11396
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 4779 10364 5087 10373
rect 4779 10362 4785 10364
rect 4841 10362 4865 10364
rect 4921 10362 4945 10364
rect 5001 10362 5025 10364
rect 5081 10362 5087 10364
rect 4841 10310 4843 10362
rect 5023 10310 5025 10362
rect 4779 10308 4785 10310
rect 4841 10308 4865 10310
rect 4921 10308 4945 10310
rect 5001 10308 5025 10310
rect 5081 10308 5087 10310
rect 4779 10299 5087 10308
rect 4779 9276 5087 9285
rect 4779 9274 4785 9276
rect 4841 9274 4865 9276
rect 4921 9274 4945 9276
rect 5001 9274 5025 9276
rect 5081 9274 5087 9276
rect 4841 9222 4843 9274
rect 5023 9222 5025 9274
rect 4779 9220 4785 9222
rect 4841 9220 4865 9222
rect 4921 9220 4945 9222
rect 5001 9220 5025 9222
rect 5081 9220 5087 9222
rect 4779 9211 5087 9220
rect 4779 8188 5087 8197
rect 4779 8186 4785 8188
rect 4841 8186 4865 8188
rect 4921 8186 4945 8188
rect 5001 8186 5025 8188
rect 5081 8186 5087 8188
rect 4841 8134 4843 8186
rect 5023 8134 5025 8186
rect 4779 8132 4785 8134
rect 4841 8132 4865 8134
rect 4921 8132 4945 8134
rect 5001 8132 5025 8134
rect 5081 8132 5087 8134
rect 4779 8123 5087 8132
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 2226 7100 2534 7109
rect 2226 7098 2232 7100
rect 2288 7098 2312 7100
rect 2368 7098 2392 7100
rect 2448 7098 2472 7100
rect 2528 7098 2534 7100
rect 2288 7046 2290 7098
rect 2470 7046 2472 7098
rect 2226 7044 2232 7046
rect 2288 7044 2312 7046
rect 2368 7044 2392 7046
rect 2448 7044 2472 7046
rect 2528 7044 2534 7046
rect 2226 7035 2534 7044
rect 4779 7100 5087 7109
rect 4779 7098 4785 7100
rect 4841 7098 4865 7100
rect 4921 7098 4945 7100
rect 5001 7098 5025 7100
rect 5081 7098 5087 7100
rect 4841 7046 4843 7098
rect 5023 7046 5025 7098
rect 4779 7044 4785 7046
rect 4841 7044 4865 7046
rect 4921 7044 4945 7046
rect 5001 7044 5025 7046
rect 5081 7044 5087 7046
rect 4779 7035 5087 7044
rect 3502 6556 3810 6565
rect 3502 6554 3508 6556
rect 3564 6554 3588 6556
rect 3644 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3810 6556
rect 3564 6502 3566 6554
rect 3746 6502 3748 6554
rect 3502 6500 3508 6502
rect 3564 6500 3588 6502
rect 3644 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3810 6502
rect 3502 6491 3810 6500
rect 2226 6012 2534 6021
rect 2226 6010 2232 6012
rect 2288 6010 2312 6012
rect 2368 6010 2392 6012
rect 2448 6010 2472 6012
rect 2528 6010 2534 6012
rect 2288 5958 2290 6010
rect 2470 5958 2472 6010
rect 2226 5956 2232 5958
rect 2288 5956 2312 5958
rect 2368 5956 2392 5958
rect 2448 5956 2472 5958
rect 2528 5956 2534 5958
rect 2226 5947 2534 5956
rect 4779 6012 5087 6021
rect 4779 6010 4785 6012
rect 4841 6010 4865 6012
rect 4921 6010 4945 6012
rect 5001 6010 5025 6012
rect 5081 6010 5087 6012
rect 4841 5958 4843 6010
rect 5023 5958 5025 6010
rect 4779 5956 4785 5958
rect 4841 5956 4865 5958
rect 4921 5956 4945 5958
rect 5001 5956 5025 5958
rect 5081 5956 5087 5958
rect 4779 5947 5087 5956
rect 3502 5468 3810 5477
rect 3502 5466 3508 5468
rect 3564 5466 3588 5468
rect 3644 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3810 5468
rect 3564 5414 3566 5466
rect 3746 5414 3748 5466
rect 3502 5412 3508 5414
rect 3564 5412 3588 5414
rect 3644 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3810 5414
rect 3502 5403 3810 5412
rect 2226 4924 2534 4933
rect 2226 4922 2232 4924
rect 2288 4922 2312 4924
rect 2368 4922 2392 4924
rect 2448 4922 2472 4924
rect 2528 4922 2534 4924
rect 2288 4870 2290 4922
rect 2470 4870 2472 4922
rect 2226 4868 2232 4870
rect 2288 4868 2312 4870
rect 2368 4868 2392 4870
rect 2448 4868 2472 4870
rect 2528 4868 2534 4870
rect 2226 4859 2534 4868
rect 4779 4924 5087 4933
rect 4779 4922 4785 4924
rect 4841 4922 4865 4924
rect 4921 4922 4945 4924
rect 5001 4922 5025 4924
rect 5081 4922 5087 4924
rect 4841 4870 4843 4922
rect 5023 4870 5025 4922
rect 4779 4868 4785 4870
rect 4841 4868 4865 4870
rect 4921 4868 4945 4870
rect 5001 4868 5025 4870
rect 5081 4868 5087 4870
rect 4779 4859 5087 4868
rect 3502 4380 3810 4389
rect 3502 4378 3508 4380
rect 3564 4378 3588 4380
rect 3644 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3810 4380
rect 3564 4326 3566 4378
rect 3746 4326 3748 4378
rect 3502 4324 3508 4326
rect 3564 4324 3588 4326
rect 3644 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3810 4326
rect 3502 4315 3810 4324
rect 2226 3836 2534 3845
rect 2226 3834 2232 3836
rect 2288 3834 2312 3836
rect 2368 3834 2392 3836
rect 2448 3834 2472 3836
rect 2528 3834 2534 3836
rect 2288 3782 2290 3834
rect 2470 3782 2472 3834
rect 2226 3780 2232 3782
rect 2288 3780 2312 3782
rect 2368 3780 2392 3782
rect 2448 3780 2472 3782
rect 2528 3780 2534 3782
rect 2226 3771 2534 3780
rect 4779 3836 5087 3845
rect 4779 3834 4785 3836
rect 4841 3834 4865 3836
rect 4921 3834 4945 3836
rect 5001 3834 5025 3836
rect 5081 3834 5087 3836
rect 4841 3782 4843 3834
rect 5023 3782 5025 3834
rect 4779 3780 4785 3782
rect 4841 3780 4865 3782
rect 4921 3780 4945 3782
rect 5001 3780 5025 3782
rect 5081 3780 5087 3782
rect 4779 3771 5087 3780
rect 5368 3738 5396 10474
rect 5552 8090 5580 10542
rect 5644 8634 5672 11018
rect 6055 10908 6363 10917
rect 6055 10906 6061 10908
rect 6117 10906 6141 10908
rect 6197 10906 6221 10908
rect 6277 10906 6301 10908
rect 6357 10906 6363 10908
rect 6117 10854 6119 10906
rect 6299 10854 6301 10906
rect 6055 10852 6061 10854
rect 6117 10852 6141 10854
rect 6197 10852 6221 10854
rect 6277 10852 6301 10854
rect 6357 10852 6363 10854
rect 6055 10843 6363 10852
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 6055 9820 6363 9829
rect 6055 9818 6061 9820
rect 6117 9818 6141 9820
rect 6197 9818 6221 9820
rect 6277 9818 6301 9820
rect 6357 9818 6363 9820
rect 6117 9766 6119 9818
rect 6299 9766 6301 9818
rect 6055 9764 6061 9766
rect 6117 9764 6141 9766
rect 6197 9764 6221 9766
rect 6277 9764 6301 9766
rect 6357 9764 6363 9766
rect 6055 9755 6363 9764
rect 6055 8732 6363 8741
rect 6055 8730 6061 8732
rect 6117 8730 6141 8732
rect 6197 8730 6221 8732
rect 6277 8730 6301 8732
rect 6357 8730 6363 8732
rect 6117 8678 6119 8730
rect 6299 8678 6301 8730
rect 6055 8676 6061 8678
rect 6117 8676 6141 8678
rect 6197 8676 6221 8678
rect 6277 8676 6301 8678
rect 6357 8676 6363 8678
rect 6055 8667 6363 8676
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 6055 7644 6363 7653
rect 6055 7642 6061 7644
rect 6117 7642 6141 7644
rect 6197 7642 6221 7644
rect 6277 7642 6301 7644
rect 6357 7642 6363 7644
rect 6117 7590 6119 7642
rect 6299 7590 6301 7642
rect 6055 7588 6061 7590
rect 6117 7588 6141 7590
rect 6197 7588 6221 7590
rect 6277 7588 6301 7590
rect 6357 7588 6363 7590
rect 6055 7579 6363 7588
rect 6055 6556 6363 6565
rect 6055 6554 6061 6556
rect 6117 6554 6141 6556
rect 6197 6554 6221 6556
rect 6277 6554 6301 6556
rect 6357 6554 6363 6556
rect 6117 6502 6119 6554
rect 6299 6502 6301 6554
rect 6055 6500 6061 6502
rect 6117 6500 6141 6502
rect 6197 6500 6221 6502
rect 6277 6500 6301 6502
rect 6357 6500 6363 6502
rect 6055 6491 6363 6500
rect 6055 5468 6363 5477
rect 6055 5466 6061 5468
rect 6117 5466 6141 5468
rect 6197 5466 6221 5468
rect 6277 5466 6301 5468
rect 6357 5466 6363 5468
rect 6117 5414 6119 5466
rect 6299 5414 6301 5466
rect 6055 5412 6061 5414
rect 6117 5412 6141 5414
rect 6197 5412 6221 5414
rect 6277 5412 6301 5414
rect 6357 5412 6363 5414
rect 6055 5403 6363 5412
rect 6055 4380 6363 4389
rect 6055 4378 6061 4380
rect 6117 4378 6141 4380
rect 6197 4378 6221 4380
rect 6277 4378 6301 4380
rect 6357 4378 6363 4380
rect 6117 4326 6119 4378
rect 6299 4326 6301 4378
rect 6055 4324 6061 4326
rect 6117 4324 6141 4326
rect 6197 4324 6221 4326
rect 6277 4324 6301 4326
rect 6357 4324 6363 4326
rect 6055 4315 6363 4324
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 1860 3664 1912 3670
rect 1860 3606 1912 3612
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3502 3292 3810 3301
rect 3502 3290 3508 3292
rect 3564 3290 3588 3292
rect 3644 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3810 3292
rect 3564 3238 3566 3290
rect 3746 3238 3748 3290
rect 3502 3236 3508 3238
rect 3564 3236 3588 3238
rect 3644 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3810 3238
rect 3502 3227 3810 3236
rect 2226 2748 2534 2757
rect 2226 2746 2232 2748
rect 2288 2746 2312 2748
rect 2368 2746 2392 2748
rect 2448 2746 2472 2748
rect 2528 2746 2534 2748
rect 2288 2694 2290 2746
rect 2470 2694 2472 2746
rect 2226 2692 2232 2694
rect 2288 2692 2312 2694
rect 2368 2692 2392 2694
rect 2448 2692 2472 2694
rect 2528 2692 2534 2694
rect 2226 2683 2534 2692
rect 4172 2650 4200 3402
rect 6055 3292 6363 3301
rect 6055 3290 6061 3292
rect 6117 3290 6141 3292
rect 6197 3290 6221 3292
rect 6277 3290 6301 3292
rect 6357 3290 6363 3292
rect 6117 3238 6119 3290
rect 6299 3238 6301 3290
rect 6055 3236 6061 3238
rect 6117 3236 6141 3238
rect 6197 3236 6221 3238
rect 6277 3236 6301 3238
rect 6357 3236 6363 3238
rect 6055 3227 6363 3236
rect 4779 2748 5087 2757
rect 4779 2746 4785 2748
rect 4841 2746 4865 2748
rect 4921 2746 4945 2748
rect 5001 2746 5025 2748
rect 5081 2746 5087 2748
rect 4841 2694 4843 2746
rect 5023 2694 5025 2746
rect 4779 2692 4785 2694
rect 4841 2692 4865 2694
rect 4921 2692 4945 2694
rect 5001 2692 5025 2694
rect 5081 2692 5087 2694
rect 4779 2683 5087 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 6564 2446 6592 8298
rect 7208 4146 7236 10746
rect 7332 10364 7640 10373
rect 7332 10362 7338 10364
rect 7394 10362 7418 10364
rect 7474 10362 7498 10364
rect 7554 10362 7578 10364
rect 7634 10362 7640 10364
rect 7394 10310 7396 10362
rect 7576 10310 7578 10362
rect 7332 10308 7338 10310
rect 7394 10308 7418 10310
rect 7474 10308 7498 10310
rect 7554 10308 7578 10310
rect 7634 10308 7640 10310
rect 7332 10299 7640 10308
rect 7332 9276 7640 9285
rect 7332 9274 7338 9276
rect 7394 9274 7418 9276
rect 7474 9274 7498 9276
rect 7554 9274 7578 9276
rect 7634 9274 7640 9276
rect 7394 9222 7396 9274
rect 7576 9222 7578 9274
rect 7332 9220 7338 9222
rect 7394 9220 7418 9222
rect 7474 9220 7498 9222
rect 7554 9220 7578 9222
rect 7634 9220 7640 9222
rect 7332 9211 7640 9220
rect 8312 9178 8340 11698
rect 9885 11452 10193 11461
rect 9885 11450 9891 11452
rect 9947 11450 9971 11452
rect 10027 11450 10051 11452
rect 10107 11450 10131 11452
rect 10187 11450 10193 11452
rect 9947 11398 9949 11450
rect 10129 11398 10131 11450
rect 9885 11396 9891 11398
rect 9947 11396 9971 11398
rect 10027 11396 10051 11398
rect 10107 11396 10131 11398
rect 10187 11396 10193 11398
rect 9885 11387 10193 11396
rect 8608 10908 8916 10917
rect 8608 10906 8614 10908
rect 8670 10906 8694 10908
rect 8750 10906 8774 10908
rect 8830 10906 8854 10908
rect 8910 10906 8916 10908
rect 8670 10854 8672 10906
rect 8852 10854 8854 10906
rect 8608 10852 8614 10854
rect 8670 10852 8694 10854
rect 8750 10852 8774 10854
rect 8830 10852 8854 10854
rect 8910 10852 8916 10854
rect 8608 10843 8916 10852
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 8608 9820 8916 9829
rect 8608 9818 8614 9820
rect 8670 9818 8694 9820
rect 8750 9818 8774 9820
rect 8830 9818 8854 9820
rect 8910 9818 8916 9820
rect 8670 9766 8672 9818
rect 8852 9766 8854 9818
rect 8608 9764 8614 9766
rect 8670 9764 8694 9766
rect 8750 9764 8774 9766
rect 8830 9764 8854 9766
rect 8910 9764 8916 9766
rect 8608 9755 8916 9764
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7332 8188 7640 8197
rect 7332 8186 7338 8188
rect 7394 8186 7418 8188
rect 7474 8186 7498 8188
rect 7554 8186 7578 8188
rect 7634 8186 7640 8188
rect 7394 8134 7396 8186
rect 7576 8134 7578 8186
rect 7332 8132 7338 8134
rect 7394 8132 7418 8134
rect 7474 8132 7498 8134
rect 7554 8132 7578 8134
rect 7634 8132 7640 8134
rect 7332 8123 7640 8132
rect 7332 7100 7640 7109
rect 7332 7098 7338 7100
rect 7394 7098 7418 7100
rect 7474 7098 7498 7100
rect 7554 7098 7578 7100
rect 7634 7098 7640 7100
rect 7394 7046 7396 7098
rect 7576 7046 7578 7098
rect 7332 7044 7338 7046
rect 7394 7044 7418 7046
rect 7474 7044 7498 7046
rect 7554 7044 7578 7046
rect 7634 7044 7640 7046
rect 7332 7035 7640 7044
rect 7332 6012 7640 6021
rect 7332 6010 7338 6012
rect 7394 6010 7418 6012
rect 7474 6010 7498 6012
rect 7554 6010 7578 6012
rect 7634 6010 7640 6012
rect 7394 5958 7396 6010
rect 7576 5958 7578 6010
rect 7332 5956 7338 5958
rect 7394 5956 7418 5958
rect 7474 5956 7498 5958
rect 7554 5956 7578 5958
rect 7634 5956 7640 5958
rect 7332 5947 7640 5956
rect 7332 4924 7640 4933
rect 7332 4922 7338 4924
rect 7394 4922 7418 4924
rect 7474 4922 7498 4924
rect 7554 4922 7578 4924
rect 7634 4922 7640 4924
rect 7394 4870 7396 4922
rect 7576 4870 7578 4922
rect 7332 4868 7338 4870
rect 7394 4868 7418 4870
rect 7474 4868 7498 4870
rect 7554 4868 7578 4870
rect 7634 4868 7640 4870
rect 7332 4859 7640 4868
rect 7668 4554 7696 8366
rect 7852 7818 7880 8434
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 7954 8248 8366
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8404 7886 8432 9318
rect 8608 8732 8916 8741
rect 8608 8730 8614 8732
rect 8670 8730 8694 8732
rect 8750 8730 8774 8732
rect 8830 8730 8854 8732
rect 8910 8730 8916 8732
rect 8670 8678 8672 8730
rect 8852 8678 8854 8730
rect 8608 8676 8614 8678
rect 8670 8676 8694 8678
rect 8750 8676 8774 8678
rect 8830 8676 8854 8678
rect 8910 8676 8916 8678
rect 8608 8667 8916 8676
rect 9324 8498 9352 10678
rect 9885 10364 10193 10373
rect 9885 10362 9891 10364
rect 9947 10362 9971 10364
rect 10027 10362 10051 10364
rect 10107 10362 10131 10364
rect 10187 10362 10193 10364
rect 9947 10310 9949 10362
rect 10129 10310 10131 10362
rect 9885 10308 9891 10310
rect 9947 10308 9971 10310
rect 10027 10308 10051 10310
rect 10107 10308 10131 10310
rect 10187 10308 10193 10310
rect 9885 10299 10193 10308
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7852 4758 7880 7754
rect 8404 7478 8432 7822
rect 8608 7644 8916 7653
rect 8608 7642 8614 7644
rect 8670 7642 8694 7644
rect 8750 7642 8774 7644
rect 8830 7642 8854 7644
rect 8910 7642 8916 7644
rect 8670 7590 8672 7642
rect 8852 7590 8854 7642
rect 8608 7588 8614 7590
rect 8670 7588 8694 7590
rect 8750 7588 8774 7590
rect 8830 7588 8854 7590
rect 8910 7588 8916 7590
rect 8608 7579 8916 7588
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 9324 6914 9352 8434
rect 9324 6886 9444 6914
rect 8608 6556 8916 6565
rect 8608 6554 8614 6556
rect 8670 6554 8694 6556
rect 8750 6554 8774 6556
rect 8830 6554 8854 6556
rect 8910 6554 8916 6556
rect 8670 6502 8672 6554
rect 8852 6502 8854 6554
rect 8608 6500 8614 6502
rect 8670 6500 8694 6502
rect 8750 6500 8774 6502
rect 8830 6500 8854 6502
rect 8910 6500 8916 6502
rect 8608 6491 8916 6500
rect 9416 5914 9444 6886
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 8608 5468 8916 5477
rect 8608 5466 8614 5468
rect 8670 5466 8694 5468
rect 8750 5466 8774 5468
rect 8830 5466 8854 5468
rect 8910 5466 8916 5468
rect 8670 5414 8672 5466
rect 8852 5414 8854 5466
rect 8608 5412 8614 5414
rect 8670 5412 8694 5414
rect 8750 5412 8774 5414
rect 8830 5412 8854 5414
rect 8910 5412 8916 5414
rect 8608 5403 8916 5412
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7332 3836 7640 3845
rect 7332 3834 7338 3836
rect 7394 3834 7418 3836
rect 7474 3834 7498 3836
rect 7554 3834 7578 3836
rect 7634 3834 7640 3836
rect 7394 3782 7396 3834
rect 7576 3782 7578 3834
rect 7332 3780 7338 3782
rect 7394 3780 7418 3782
rect 7474 3780 7498 3782
rect 7554 3780 7578 3782
rect 7634 3780 7640 3782
rect 7332 3771 7640 3780
rect 7668 3466 7696 4490
rect 7852 3602 7880 4694
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 8608 4380 8916 4389
rect 8608 4378 8614 4380
rect 8670 4378 8694 4380
rect 8750 4378 8774 4380
rect 8830 4378 8854 4380
rect 8910 4378 8916 4380
rect 8670 4326 8672 4378
rect 8852 4326 8854 4378
rect 8608 4324 8614 4326
rect 8670 4324 8694 4326
rect 8750 4324 8774 4326
rect 8830 4324 8854 4326
rect 8910 4324 8916 4326
rect 8608 4315 8916 4324
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 9324 3534 9352 4422
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 8608 3292 8916 3301
rect 8608 3290 8614 3292
rect 8670 3290 8694 3292
rect 8750 3290 8774 3292
rect 8830 3290 8854 3292
rect 8910 3290 8916 3292
rect 8670 3238 8672 3290
rect 8852 3238 8854 3290
rect 8608 3236 8614 3238
rect 8670 3236 8694 3238
rect 8750 3236 8774 3238
rect 8830 3236 8854 3238
rect 8910 3236 8916 3238
rect 8608 3227 8916 3236
rect 9692 3058 9720 9522
rect 9885 9276 10193 9285
rect 9885 9274 9891 9276
rect 9947 9274 9971 9276
rect 10027 9274 10051 9276
rect 10107 9274 10131 9276
rect 10187 9274 10193 9276
rect 9947 9222 9949 9274
rect 10129 9222 10131 9274
rect 9885 9220 9891 9222
rect 9947 9220 9971 9222
rect 10027 9220 10051 9222
rect 10107 9220 10131 9222
rect 10187 9220 10193 9222
rect 9885 9211 10193 9220
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 9885 8188 10193 8197
rect 9885 8186 9891 8188
rect 9947 8186 9971 8188
rect 10027 8186 10051 8188
rect 10107 8186 10131 8188
rect 10187 8186 10193 8188
rect 9947 8134 9949 8186
rect 10129 8134 10131 8186
rect 9885 8132 9891 8134
rect 9947 8132 9971 8134
rect 10027 8132 10051 8134
rect 10107 8132 10131 8134
rect 10187 8132 10193 8134
rect 9885 8123 10193 8132
rect 10428 8090 10456 8366
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9784 3738 9812 7346
rect 9885 7100 10193 7109
rect 9885 7098 9891 7100
rect 9947 7098 9971 7100
rect 10027 7098 10051 7100
rect 10107 7098 10131 7100
rect 10187 7098 10193 7100
rect 9947 7046 9949 7098
rect 10129 7046 10131 7098
rect 9885 7044 9891 7046
rect 9947 7044 9971 7046
rect 10027 7044 10051 7046
rect 10107 7044 10131 7046
rect 10187 7044 10193 7046
rect 9885 7035 10193 7044
rect 9885 6012 10193 6021
rect 9885 6010 9891 6012
rect 9947 6010 9971 6012
rect 10027 6010 10051 6012
rect 10107 6010 10131 6012
rect 10187 6010 10193 6012
rect 9947 5958 9949 6010
rect 10129 5958 10131 6010
rect 9885 5956 9891 5958
rect 9947 5956 9971 5958
rect 10027 5956 10051 5958
rect 10107 5956 10131 5958
rect 10187 5956 10193 5958
rect 9885 5947 10193 5956
rect 9885 4924 10193 4933
rect 9885 4922 9891 4924
rect 9947 4922 9971 4924
rect 10027 4922 10051 4924
rect 10107 4922 10131 4924
rect 10187 4922 10193 4924
rect 9947 4870 9949 4922
rect 10129 4870 10131 4922
rect 9885 4868 9891 4870
rect 9947 4868 9971 4870
rect 10027 4868 10051 4870
rect 10107 4868 10131 4870
rect 10187 4868 10193 4870
rect 9885 4859 10193 4868
rect 10520 4010 10548 11698
rect 10690 11656 10746 11665
rect 10690 11591 10692 11600
rect 10744 11591 10746 11600
rect 10692 11562 10744 11568
rect 11161 10908 11469 10917
rect 11161 10906 11167 10908
rect 11223 10906 11247 10908
rect 11303 10906 11327 10908
rect 11383 10906 11407 10908
rect 11463 10906 11469 10908
rect 11223 10854 11225 10906
rect 11405 10854 11407 10906
rect 11161 10852 11167 10854
rect 11223 10852 11247 10854
rect 11303 10852 11327 10854
rect 11383 10852 11407 10854
rect 11463 10852 11469 10854
rect 11161 10843 11469 10852
rect 11161 9820 11469 9829
rect 11161 9818 11167 9820
rect 11223 9818 11247 9820
rect 11303 9818 11327 9820
rect 11383 9818 11407 9820
rect 11463 9818 11469 9820
rect 11223 9766 11225 9818
rect 11405 9766 11407 9818
rect 11161 9764 11167 9766
rect 11223 9764 11247 9766
rect 11303 9764 11327 9766
rect 11383 9764 11407 9766
rect 11463 9764 11469 9766
rect 11161 9755 11469 9764
rect 11161 8732 11469 8741
rect 11161 8730 11167 8732
rect 11223 8730 11247 8732
rect 11303 8730 11327 8732
rect 11383 8730 11407 8732
rect 11463 8730 11469 8732
rect 11223 8678 11225 8730
rect 11405 8678 11407 8730
rect 11161 8676 11167 8678
rect 11223 8676 11247 8678
rect 11303 8676 11327 8678
rect 11383 8676 11407 8678
rect 11463 8676 11469 8678
rect 11161 8667 11469 8676
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 7478 10732 8366
rect 11161 7644 11469 7653
rect 11161 7642 11167 7644
rect 11223 7642 11247 7644
rect 11303 7642 11327 7644
rect 11383 7642 11407 7644
rect 11463 7642 11469 7644
rect 11223 7590 11225 7642
rect 11405 7590 11407 7642
rect 11161 7588 11167 7590
rect 11223 7588 11247 7590
rect 11303 7588 11327 7590
rect 11383 7588 11407 7590
rect 11463 7588 11469 7590
rect 11161 7579 11469 7588
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 11161 6556 11469 6565
rect 11161 6554 11167 6556
rect 11223 6554 11247 6556
rect 11303 6554 11327 6556
rect 11383 6554 11407 6556
rect 11463 6554 11469 6556
rect 11223 6502 11225 6554
rect 11405 6502 11407 6554
rect 11161 6500 11167 6502
rect 11223 6500 11247 6502
rect 11303 6500 11327 6502
rect 11383 6500 11407 6502
rect 11463 6500 11469 6502
rect 11161 6491 11469 6500
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5273 10824 5646
rect 11161 5468 11469 5477
rect 11161 5466 11167 5468
rect 11223 5466 11247 5468
rect 11303 5466 11327 5468
rect 11383 5466 11407 5468
rect 11463 5466 11469 5468
rect 11223 5414 11225 5466
rect 11405 5414 11407 5466
rect 11161 5412 11167 5414
rect 11223 5412 11247 5414
rect 11303 5412 11327 5414
rect 11383 5412 11407 5414
rect 11463 5412 11469 5414
rect 11161 5403 11469 5412
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 11161 4380 11469 4389
rect 11161 4378 11167 4380
rect 11223 4378 11247 4380
rect 11303 4378 11327 4380
rect 11383 4378 11407 4380
rect 11463 4378 11469 4380
rect 11223 4326 11225 4378
rect 11405 4326 11407 4378
rect 11161 4324 11167 4326
rect 11223 4324 11247 4326
rect 11303 4324 11327 4326
rect 11383 4324 11407 4326
rect 11463 4324 11469 4326
rect 11161 4315 11469 4324
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 9885 3836 10193 3845
rect 9885 3834 9891 3836
rect 9947 3834 9971 3836
rect 10027 3834 10051 3836
rect 10107 3834 10131 3836
rect 10187 3834 10193 3836
rect 9947 3782 9949 3834
rect 10129 3782 10131 3834
rect 9885 3780 9891 3782
rect 9947 3780 9971 3782
rect 10027 3780 10051 3782
rect 10107 3780 10131 3782
rect 10187 3780 10193 3782
rect 9885 3771 10193 3780
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 11161 3292 11469 3301
rect 11161 3290 11167 3292
rect 11223 3290 11247 3292
rect 11303 3290 11327 3292
rect 11383 3290 11407 3292
rect 11463 3290 11469 3292
rect 11223 3238 11225 3290
rect 11405 3238 11407 3290
rect 11161 3236 11167 3238
rect 11223 3236 11247 3238
rect 11303 3236 11327 3238
rect 11383 3236 11407 3238
rect 11463 3236 11469 3238
rect 11161 3227 11469 3236
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 7332 2748 7640 2757
rect 7332 2746 7338 2748
rect 7394 2746 7418 2748
rect 7474 2746 7498 2748
rect 7554 2746 7578 2748
rect 7634 2746 7640 2748
rect 7394 2694 7396 2746
rect 7576 2694 7578 2746
rect 7332 2692 7338 2694
rect 7394 2692 7418 2694
rect 7474 2692 7498 2694
rect 7554 2692 7578 2694
rect 7634 2692 7640 2694
rect 7332 2683 7640 2692
rect 9885 2748 10193 2757
rect 9885 2746 9891 2748
rect 9947 2746 9971 2748
rect 10027 2746 10051 2748
rect 10107 2746 10131 2748
rect 10187 2746 10193 2748
rect 9947 2694 9949 2746
rect 10129 2694 10131 2746
rect 9885 2692 9891 2694
rect 9947 2692 9971 2694
rect 10027 2692 10051 2694
rect 10107 2692 10131 2694
rect 10187 2692 10193 2694
rect 9885 2683 10193 2692
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 32 800 60 2382
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 3502 2204 3810 2213
rect 3502 2202 3508 2204
rect 3564 2202 3588 2204
rect 3644 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3810 2204
rect 3564 2150 3566 2202
rect 3746 2150 3748 2202
rect 3502 2148 3508 2150
rect 3564 2148 3588 2150
rect 3644 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3810 2150
rect 3502 2139 3810 2148
rect 5828 800 5856 2246
rect 6055 2204 6363 2213
rect 6055 2202 6061 2204
rect 6117 2202 6141 2204
rect 6197 2202 6221 2204
rect 6277 2202 6301 2204
rect 6357 2202 6363 2204
rect 6117 2150 6119 2202
rect 6299 2150 6301 2202
rect 6055 2148 6061 2150
rect 6117 2148 6141 2150
rect 6197 2148 6221 2150
rect 6277 2148 6301 2150
rect 6357 2148 6363 2150
rect 6055 2139 6363 2148
rect 8608 2204 8916 2213
rect 8608 2202 8614 2204
rect 8670 2202 8694 2204
rect 8750 2202 8774 2204
rect 8830 2202 8854 2204
rect 8910 2202 8916 2204
rect 8670 2150 8672 2202
rect 8852 2150 8854 2202
rect 8608 2148 8614 2150
rect 8670 2148 8694 2150
rect 8750 2148 8774 2150
rect 8830 2148 8854 2150
rect 8910 2148 8916 2150
rect 8608 2139 8916 2148
rect 11161 2204 11469 2213
rect 11161 2202 11167 2204
rect 11223 2202 11247 2204
rect 11303 2202 11327 2204
rect 11383 2202 11407 2204
rect 11463 2202 11469 2204
rect 11223 2150 11225 2202
rect 11405 2150 11407 2202
rect 11161 2148 11167 2150
rect 11223 2148 11247 2150
rect 11303 2148 11327 2150
rect 11383 2148 11407 2150
rect 11463 2148 11469 2150
rect 11161 2139 11469 2148
rect 11624 800 11652 2994
rect 18 0 74 800
rect 5814 0 5870 800
rect 11610 0 11666 800
<< via2 >>
rect 1674 12280 1730 12336
rect 3508 11994 3564 11996
rect 3588 11994 3644 11996
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3508 11942 3554 11994
rect 3554 11942 3564 11994
rect 3588 11942 3618 11994
rect 3618 11942 3630 11994
rect 3630 11942 3644 11994
rect 3668 11942 3682 11994
rect 3682 11942 3694 11994
rect 3694 11942 3724 11994
rect 3748 11942 3758 11994
rect 3758 11942 3804 11994
rect 3508 11940 3564 11942
rect 3588 11940 3644 11942
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 6061 11994 6117 11996
rect 6141 11994 6197 11996
rect 6221 11994 6277 11996
rect 6301 11994 6357 11996
rect 6061 11942 6107 11994
rect 6107 11942 6117 11994
rect 6141 11942 6171 11994
rect 6171 11942 6183 11994
rect 6183 11942 6197 11994
rect 6221 11942 6235 11994
rect 6235 11942 6247 11994
rect 6247 11942 6277 11994
rect 6301 11942 6311 11994
rect 6311 11942 6357 11994
rect 6061 11940 6117 11942
rect 6141 11940 6197 11942
rect 6221 11940 6277 11942
rect 6301 11940 6357 11942
rect 8614 11994 8670 11996
rect 8694 11994 8750 11996
rect 8774 11994 8830 11996
rect 8854 11994 8910 11996
rect 8614 11942 8660 11994
rect 8660 11942 8670 11994
rect 8694 11942 8724 11994
rect 8724 11942 8736 11994
rect 8736 11942 8750 11994
rect 8774 11942 8788 11994
rect 8788 11942 8800 11994
rect 8800 11942 8830 11994
rect 8854 11942 8864 11994
rect 8864 11942 8910 11994
rect 8614 11940 8670 11942
rect 8694 11940 8750 11942
rect 8774 11940 8830 11942
rect 8854 11940 8910 11942
rect 11167 11994 11223 11996
rect 11247 11994 11303 11996
rect 11327 11994 11383 11996
rect 11407 11994 11463 11996
rect 11167 11942 11213 11994
rect 11213 11942 11223 11994
rect 11247 11942 11277 11994
rect 11277 11942 11289 11994
rect 11289 11942 11303 11994
rect 11327 11942 11341 11994
rect 11341 11942 11353 11994
rect 11353 11942 11383 11994
rect 11407 11942 11417 11994
rect 11417 11942 11463 11994
rect 11167 11940 11223 11942
rect 11247 11940 11303 11942
rect 11327 11940 11383 11942
rect 11407 11940 11463 11942
rect 2232 11450 2288 11452
rect 2312 11450 2368 11452
rect 2392 11450 2448 11452
rect 2472 11450 2528 11452
rect 2232 11398 2278 11450
rect 2278 11398 2288 11450
rect 2312 11398 2342 11450
rect 2342 11398 2354 11450
rect 2354 11398 2368 11450
rect 2392 11398 2406 11450
rect 2406 11398 2418 11450
rect 2418 11398 2448 11450
rect 2472 11398 2482 11450
rect 2482 11398 2528 11450
rect 2232 11396 2288 11398
rect 2312 11396 2368 11398
rect 2392 11396 2448 11398
rect 2472 11396 2528 11398
rect 3508 10906 3564 10908
rect 3588 10906 3644 10908
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3508 10854 3554 10906
rect 3554 10854 3564 10906
rect 3588 10854 3618 10906
rect 3618 10854 3630 10906
rect 3630 10854 3644 10906
rect 3668 10854 3682 10906
rect 3682 10854 3694 10906
rect 3694 10854 3724 10906
rect 3748 10854 3758 10906
rect 3758 10854 3804 10906
rect 3508 10852 3564 10854
rect 3588 10852 3644 10854
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 2232 10362 2288 10364
rect 2312 10362 2368 10364
rect 2392 10362 2448 10364
rect 2472 10362 2528 10364
rect 2232 10310 2278 10362
rect 2278 10310 2288 10362
rect 2312 10310 2342 10362
rect 2342 10310 2354 10362
rect 2354 10310 2368 10362
rect 2392 10310 2406 10362
rect 2406 10310 2418 10362
rect 2418 10310 2448 10362
rect 2472 10310 2482 10362
rect 2482 10310 2528 10362
rect 2232 10308 2288 10310
rect 2312 10308 2368 10310
rect 2392 10308 2448 10310
rect 2472 10308 2528 10310
rect 3508 9818 3564 9820
rect 3588 9818 3644 9820
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3508 9766 3554 9818
rect 3554 9766 3564 9818
rect 3588 9766 3618 9818
rect 3618 9766 3630 9818
rect 3630 9766 3644 9818
rect 3668 9766 3682 9818
rect 3682 9766 3694 9818
rect 3694 9766 3724 9818
rect 3748 9766 3758 9818
rect 3758 9766 3804 9818
rect 3508 9764 3564 9766
rect 3588 9764 3644 9766
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 2232 9274 2288 9276
rect 2312 9274 2368 9276
rect 2392 9274 2448 9276
rect 2472 9274 2528 9276
rect 2232 9222 2278 9274
rect 2278 9222 2288 9274
rect 2312 9222 2342 9274
rect 2342 9222 2354 9274
rect 2354 9222 2368 9274
rect 2392 9222 2406 9274
rect 2406 9222 2418 9274
rect 2418 9222 2448 9274
rect 2472 9222 2482 9274
rect 2482 9222 2528 9274
rect 2232 9220 2288 9222
rect 2312 9220 2368 9222
rect 2392 9220 2448 9222
rect 2472 9220 2528 9222
rect 3508 8730 3564 8732
rect 3588 8730 3644 8732
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3508 8678 3554 8730
rect 3554 8678 3564 8730
rect 3588 8678 3618 8730
rect 3618 8678 3630 8730
rect 3630 8678 3644 8730
rect 3668 8678 3682 8730
rect 3682 8678 3694 8730
rect 3694 8678 3724 8730
rect 3748 8678 3758 8730
rect 3758 8678 3804 8730
rect 3508 8676 3564 8678
rect 3588 8676 3644 8678
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 2232 8186 2288 8188
rect 2312 8186 2368 8188
rect 2392 8186 2448 8188
rect 2472 8186 2528 8188
rect 2232 8134 2278 8186
rect 2278 8134 2288 8186
rect 2312 8134 2342 8186
rect 2342 8134 2354 8186
rect 2354 8134 2368 8186
rect 2392 8134 2406 8186
rect 2406 8134 2418 8186
rect 2418 8134 2448 8186
rect 2472 8134 2482 8186
rect 2482 8134 2528 8186
rect 2232 8132 2288 8134
rect 2312 8132 2368 8134
rect 2392 8132 2448 8134
rect 2472 8132 2528 8134
rect 3508 7642 3564 7644
rect 3588 7642 3644 7644
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3508 7590 3554 7642
rect 3554 7590 3564 7642
rect 3588 7590 3618 7642
rect 3618 7590 3630 7642
rect 3630 7590 3644 7642
rect 3668 7590 3682 7642
rect 3682 7590 3694 7642
rect 3694 7590 3724 7642
rect 3748 7590 3758 7642
rect 3758 7590 3804 7642
rect 3508 7588 3564 7590
rect 3588 7588 3644 7590
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 4785 11450 4841 11452
rect 4865 11450 4921 11452
rect 4945 11450 5001 11452
rect 5025 11450 5081 11452
rect 4785 11398 4831 11450
rect 4831 11398 4841 11450
rect 4865 11398 4895 11450
rect 4895 11398 4907 11450
rect 4907 11398 4921 11450
rect 4945 11398 4959 11450
rect 4959 11398 4971 11450
rect 4971 11398 5001 11450
rect 5025 11398 5035 11450
rect 5035 11398 5081 11450
rect 4785 11396 4841 11398
rect 4865 11396 4921 11398
rect 4945 11396 5001 11398
rect 5025 11396 5081 11398
rect 7338 11450 7394 11452
rect 7418 11450 7474 11452
rect 7498 11450 7554 11452
rect 7578 11450 7634 11452
rect 7338 11398 7384 11450
rect 7384 11398 7394 11450
rect 7418 11398 7448 11450
rect 7448 11398 7460 11450
rect 7460 11398 7474 11450
rect 7498 11398 7512 11450
rect 7512 11398 7524 11450
rect 7524 11398 7554 11450
rect 7578 11398 7588 11450
rect 7588 11398 7634 11450
rect 7338 11396 7394 11398
rect 7418 11396 7474 11398
rect 7498 11396 7554 11398
rect 7578 11396 7634 11398
rect 4785 10362 4841 10364
rect 4865 10362 4921 10364
rect 4945 10362 5001 10364
rect 5025 10362 5081 10364
rect 4785 10310 4831 10362
rect 4831 10310 4841 10362
rect 4865 10310 4895 10362
rect 4895 10310 4907 10362
rect 4907 10310 4921 10362
rect 4945 10310 4959 10362
rect 4959 10310 4971 10362
rect 4971 10310 5001 10362
rect 5025 10310 5035 10362
rect 5035 10310 5081 10362
rect 4785 10308 4841 10310
rect 4865 10308 4921 10310
rect 4945 10308 5001 10310
rect 5025 10308 5081 10310
rect 4785 9274 4841 9276
rect 4865 9274 4921 9276
rect 4945 9274 5001 9276
rect 5025 9274 5081 9276
rect 4785 9222 4831 9274
rect 4831 9222 4841 9274
rect 4865 9222 4895 9274
rect 4895 9222 4907 9274
rect 4907 9222 4921 9274
rect 4945 9222 4959 9274
rect 4959 9222 4971 9274
rect 4971 9222 5001 9274
rect 5025 9222 5035 9274
rect 5035 9222 5081 9274
rect 4785 9220 4841 9222
rect 4865 9220 4921 9222
rect 4945 9220 5001 9222
rect 5025 9220 5081 9222
rect 4785 8186 4841 8188
rect 4865 8186 4921 8188
rect 4945 8186 5001 8188
rect 5025 8186 5081 8188
rect 4785 8134 4831 8186
rect 4831 8134 4841 8186
rect 4865 8134 4895 8186
rect 4895 8134 4907 8186
rect 4907 8134 4921 8186
rect 4945 8134 4959 8186
rect 4959 8134 4971 8186
rect 4971 8134 5001 8186
rect 5025 8134 5035 8186
rect 5035 8134 5081 8186
rect 4785 8132 4841 8134
rect 4865 8132 4921 8134
rect 4945 8132 5001 8134
rect 5025 8132 5081 8134
rect 2232 7098 2288 7100
rect 2312 7098 2368 7100
rect 2392 7098 2448 7100
rect 2472 7098 2528 7100
rect 2232 7046 2278 7098
rect 2278 7046 2288 7098
rect 2312 7046 2342 7098
rect 2342 7046 2354 7098
rect 2354 7046 2368 7098
rect 2392 7046 2406 7098
rect 2406 7046 2418 7098
rect 2418 7046 2448 7098
rect 2472 7046 2482 7098
rect 2482 7046 2528 7098
rect 2232 7044 2288 7046
rect 2312 7044 2368 7046
rect 2392 7044 2448 7046
rect 2472 7044 2528 7046
rect 4785 7098 4841 7100
rect 4865 7098 4921 7100
rect 4945 7098 5001 7100
rect 5025 7098 5081 7100
rect 4785 7046 4831 7098
rect 4831 7046 4841 7098
rect 4865 7046 4895 7098
rect 4895 7046 4907 7098
rect 4907 7046 4921 7098
rect 4945 7046 4959 7098
rect 4959 7046 4971 7098
rect 4971 7046 5001 7098
rect 5025 7046 5035 7098
rect 5035 7046 5081 7098
rect 4785 7044 4841 7046
rect 4865 7044 4921 7046
rect 4945 7044 5001 7046
rect 5025 7044 5081 7046
rect 3508 6554 3564 6556
rect 3588 6554 3644 6556
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3508 6502 3554 6554
rect 3554 6502 3564 6554
rect 3588 6502 3618 6554
rect 3618 6502 3630 6554
rect 3630 6502 3644 6554
rect 3668 6502 3682 6554
rect 3682 6502 3694 6554
rect 3694 6502 3724 6554
rect 3748 6502 3758 6554
rect 3758 6502 3804 6554
rect 3508 6500 3564 6502
rect 3588 6500 3644 6502
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 2232 6010 2288 6012
rect 2312 6010 2368 6012
rect 2392 6010 2448 6012
rect 2472 6010 2528 6012
rect 2232 5958 2278 6010
rect 2278 5958 2288 6010
rect 2312 5958 2342 6010
rect 2342 5958 2354 6010
rect 2354 5958 2368 6010
rect 2392 5958 2406 6010
rect 2406 5958 2418 6010
rect 2418 5958 2448 6010
rect 2472 5958 2482 6010
rect 2482 5958 2528 6010
rect 2232 5956 2288 5958
rect 2312 5956 2368 5958
rect 2392 5956 2448 5958
rect 2472 5956 2528 5958
rect 4785 6010 4841 6012
rect 4865 6010 4921 6012
rect 4945 6010 5001 6012
rect 5025 6010 5081 6012
rect 4785 5958 4831 6010
rect 4831 5958 4841 6010
rect 4865 5958 4895 6010
rect 4895 5958 4907 6010
rect 4907 5958 4921 6010
rect 4945 5958 4959 6010
rect 4959 5958 4971 6010
rect 4971 5958 5001 6010
rect 5025 5958 5035 6010
rect 5035 5958 5081 6010
rect 4785 5956 4841 5958
rect 4865 5956 4921 5958
rect 4945 5956 5001 5958
rect 5025 5956 5081 5958
rect 3508 5466 3564 5468
rect 3588 5466 3644 5468
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3508 5414 3554 5466
rect 3554 5414 3564 5466
rect 3588 5414 3618 5466
rect 3618 5414 3630 5466
rect 3630 5414 3644 5466
rect 3668 5414 3682 5466
rect 3682 5414 3694 5466
rect 3694 5414 3724 5466
rect 3748 5414 3758 5466
rect 3758 5414 3804 5466
rect 3508 5412 3564 5414
rect 3588 5412 3644 5414
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 2232 4922 2288 4924
rect 2312 4922 2368 4924
rect 2392 4922 2448 4924
rect 2472 4922 2528 4924
rect 2232 4870 2278 4922
rect 2278 4870 2288 4922
rect 2312 4870 2342 4922
rect 2342 4870 2354 4922
rect 2354 4870 2368 4922
rect 2392 4870 2406 4922
rect 2406 4870 2418 4922
rect 2418 4870 2448 4922
rect 2472 4870 2482 4922
rect 2482 4870 2528 4922
rect 2232 4868 2288 4870
rect 2312 4868 2368 4870
rect 2392 4868 2448 4870
rect 2472 4868 2528 4870
rect 4785 4922 4841 4924
rect 4865 4922 4921 4924
rect 4945 4922 5001 4924
rect 5025 4922 5081 4924
rect 4785 4870 4831 4922
rect 4831 4870 4841 4922
rect 4865 4870 4895 4922
rect 4895 4870 4907 4922
rect 4907 4870 4921 4922
rect 4945 4870 4959 4922
rect 4959 4870 4971 4922
rect 4971 4870 5001 4922
rect 5025 4870 5035 4922
rect 5035 4870 5081 4922
rect 4785 4868 4841 4870
rect 4865 4868 4921 4870
rect 4945 4868 5001 4870
rect 5025 4868 5081 4870
rect 3508 4378 3564 4380
rect 3588 4378 3644 4380
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3508 4326 3554 4378
rect 3554 4326 3564 4378
rect 3588 4326 3618 4378
rect 3618 4326 3630 4378
rect 3630 4326 3644 4378
rect 3668 4326 3682 4378
rect 3682 4326 3694 4378
rect 3694 4326 3724 4378
rect 3748 4326 3758 4378
rect 3758 4326 3804 4378
rect 3508 4324 3564 4326
rect 3588 4324 3644 4326
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 2232 3834 2288 3836
rect 2312 3834 2368 3836
rect 2392 3834 2448 3836
rect 2472 3834 2528 3836
rect 2232 3782 2278 3834
rect 2278 3782 2288 3834
rect 2312 3782 2342 3834
rect 2342 3782 2354 3834
rect 2354 3782 2368 3834
rect 2392 3782 2406 3834
rect 2406 3782 2418 3834
rect 2418 3782 2448 3834
rect 2472 3782 2482 3834
rect 2482 3782 2528 3834
rect 2232 3780 2288 3782
rect 2312 3780 2368 3782
rect 2392 3780 2448 3782
rect 2472 3780 2528 3782
rect 4785 3834 4841 3836
rect 4865 3834 4921 3836
rect 4945 3834 5001 3836
rect 5025 3834 5081 3836
rect 4785 3782 4831 3834
rect 4831 3782 4841 3834
rect 4865 3782 4895 3834
rect 4895 3782 4907 3834
rect 4907 3782 4921 3834
rect 4945 3782 4959 3834
rect 4959 3782 4971 3834
rect 4971 3782 5001 3834
rect 5025 3782 5035 3834
rect 5035 3782 5081 3834
rect 4785 3780 4841 3782
rect 4865 3780 4921 3782
rect 4945 3780 5001 3782
rect 5025 3780 5081 3782
rect 6061 10906 6117 10908
rect 6141 10906 6197 10908
rect 6221 10906 6277 10908
rect 6301 10906 6357 10908
rect 6061 10854 6107 10906
rect 6107 10854 6117 10906
rect 6141 10854 6171 10906
rect 6171 10854 6183 10906
rect 6183 10854 6197 10906
rect 6221 10854 6235 10906
rect 6235 10854 6247 10906
rect 6247 10854 6277 10906
rect 6301 10854 6311 10906
rect 6311 10854 6357 10906
rect 6061 10852 6117 10854
rect 6141 10852 6197 10854
rect 6221 10852 6277 10854
rect 6301 10852 6357 10854
rect 6061 9818 6117 9820
rect 6141 9818 6197 9820
rect 6221 9818 6277 9820
rect 6301 9818 6357 9820
rect 6061 9766 6107 9818
rect 6107 9766 6117 9818
rect 6141 9766 6171 9818
rect 6171 9766 6183 9818
rect 6183 9766 6197 9818
rect 6221 9766 6235 9818
rect 6235 9766 6247 9818
rect 6247 9766 6277 9818
rect 6301 9766 6311 9818
rect 6311 9766 6357 9818
rect 6061 9764 6117 9766
rect 6141 9764 6197 9766
rect 6221 9764 6277 9766
rect 6301 9764 6357 9766
rect 6061 8730 6117 8732
rect 6141 8730 6197 8732
rect 6221 8730 6277 8732
rect 6301 8730 6357 8732
rect 6061 8678 6107 8730
rect 6107 8678 6117 8730
rect 6141 8678 6171 8730
rect 6171 8678 6183 8730
rect 6183 8678 6197 8730
rect 6221 8678 6235 8730
rect 6235 8678 6247 8730
rect 6247 8678 6277 8730
rect 6301 8678 6311 8730
rect 6311 8678 6357 8730
rect 6061 8676 6117 8678
rect 6141 8676 6197 8678
rect 6221 8676 6277 8678
rect 6301 8676 6357 8678
rect 6061 7642 6117 7644
rect 6141 7642 6197 7644
rect 6221 7642 6277 7644
rect 6301 7642 6357 7644
rect 6061 7590 6107 7642
rect 6107 7590 6117 7642
rect 6141 7590 6171 7642
rect 6171 7590 6183 7642
rect 6183 7590 6197 7642
rect 6221 7590 6235 7642
rect 6235 7590 6247 7642
rect 6247 7590 6277 7642
rect 6301 7590 6311 7642
rect 6311 7590 6357 7642
rect 6061 7588 6117 7590
rect 6141 7588 6197 7590
rect 6221 7588 6277 7590
rect 6301 7588 6357 7590
rect 6061 6554 6117 6556
rect 6141 6554 6197 6556
rect 6221 6554 6277 6556
rect 6301 6554 6357 6556
rect 6061 6502 6107 6554
rect 6107 6502 6117 6554
rect 6141 6502 6171 6554
rect 6171 6502 6183 6554
rect 6183 6502 6197 6554
rect 6221 6502 6235 6554
rect 6235 6502 6247 6554
rect 6247 6502 6277 6554
rect 6301 6502 6311 6554
rect 6311 6502 6357 6554
rect 6061 6500 6117 6502
rect 6141 6500 6197 6502
rect 6221 6500 6277 6502
rect 6301 6500 6357 6502
rect 6061 5466 6117 5468
rect 6141 5466 6197 5468
rect 6221 5466 6277 5468
rect 6301 5466 6357 5468
rect 6061 5414 6107 5466
rect 6107 5414 6117 5466
rect 6141 5414 6171 5466
rect 6171 5414 6183 5466
rect 6183 5414 6197 5466
rect 6221 5414 6235 5466
rect 6235 5414 6247 5466
rect 6247 5414 6277 5466
rect 6301 5414 6311 5466
rect 6311 5414 6357 5466
rect 6061 5412 6117 5414
rect 6141 5412 6197 5414
rect 6221 5412 6277 5414
rect 6301 5412 6357 5414
rect 6061 4378 6117 4380
rect 6141 4378 6197 4380
rect 6221 4378 6277 4380
rect 6301 4378 6357 4380
rect 6061 4326 6107 4378
rect 6107 4326 6117 4378
rect 6141 4326 6171 4378
rect 6171 4326 6183 4378
rect 6183 4326 6197 4378
rect 6221 4326 6235 4378
rect 6235 4326 6247 4378
rect 6247 4326 6277 4378
rect 6301 4326 6311 4378
rect 6311 4326 6357 4378
rect 6061 4324 6117 4326
rect 6141 4324 6197 4326
rect 6221 4324 6277 4326
rect 6301 4324 6357 4326
rect 3508 3290 3564 3292
rect 3588 3290 3644 3292
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3508 3238 3554 3290
rect 3554 3238 3564 3290
rect 3588 3238 3618 3290
rect 3618 3238 3630 3290
rect 3630 3238 3644 3290
rect 3668 3238 3682 3290
rect 3682 3238 3694 3290
rect 3694 3238 3724 3290
rect 3748 3238 3758 3290
rect 3758 3238 3804 3290
rect 3508 3236 3564 3238
rect 3588 3236 3644 3238
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 2232 2746 2288 2748
rect 2312 2746 2368 2748
rect 2392 2746 2448 2748
rect 2472 2746 2528 2748
rect 2232 2694 2278 2746
rect 2278 2694 2288 2746
rect 2312 2694 2342 2746
rect 2342 2694 2354 2746
rect 2354 2694 2368 2746
rect 2392 2694 2406 2746
rect 2406 2694 2418 2746
rect 2418 2694 2448 2746
rect 2472 2694 2482 2746
rect 2482 2694 2528 2746
rect 2232 2692 2288 2694
rect 2312 2692 2368 2694
rect 2392 2692 2448 2694
rect 2472 2692 2528 2694
rect 6061 3290 6117 3292
rect 6141 3290 6197 3292
rect 6221 3290 6277 3292
rect 6301 3290 6357 3292
rect 6061 3238 6107 3290
rect 6107 3238 6117 3290
rect 6141 3238 6171 3290
rect 6171 3238 6183 3290
rect 6183 3238 6197 3290
rect 6221 3238 6235 3290
rect 6235 3238 6247 3290
rect 6247 3238 6277 3290
rect 6301 3238 6311 3290
rect 6311 3238 6357 3290
rect 6061 3236 6117 3238
rect 6141 3236 6197 3238
rect 6221 3236 6277 3238
rect 6301 3236 6357 3238
rect 4785 2746 4841 2748
rect 4865 2746 4921 2748
rect 4945 2746 5001 2748
rect 5025 2746 5081 2748
rect 4785 2694 4831 2746
rect 4831 2694 4841 2746
rect 4865 2694 4895 2746
rect 4895 2694 4907 2746
rect 4907 2694 4921 2746
rect 4945 2694 4959 2746
rect 4959 2694 4971 2746
rect 4971 2694 5001 2746
rect 5025 2694 5035 2746
rect 5035 2694 5081 2746
rect 4785 2692 4841 2694
rect 4865 2692 4921 2694
rect 4945 2692 5001 2694
rect 5025 2692 5081 2694
rect 7338 10362 7394 10364
rect 7418 10362 7474 10364
rect 7498 10362 7554 10364
rect 7578 10362 7634 10364
rect 7338 10310 7384 10362
rect 7384 10310 7394 10362
rect 7418 10310 7448 10362
rect 7448 10310 7460 10362
rect 7460 10310 7474 10362
rect 7498 10310 7512 10362
rect 7512 10310 7524 10362
rect 7524 10310 7554 10362
rect 7578 10310 7588 10362
rect 7588 10310 7634 10362
rect 7338 10308 7394 10310
rect 7418 10308 7474 10310
rect 7498 10308 7554 10310
rect 7578 10308 7634 10310
rect 7338 9274 7394 9276
rect 7418 9274 7474 9276
rect 7498 9274 7554 9276
rect 7578 9274 7634 9276
rect 7338 9222 7384 9274
rect 7384 9222 7394 9274
rect 7418 9222 7448 9274
rect 7448 9222 7460 9274
rect 7460 9222 7474 9274
rect 7498 9222 7512 9274
rect 7512 9222 7524 9274
rect 7524 9222 7554 9274
rect 7578 9222 7588 9274
rect 7588 9222 7634 9274
rect 7338 9220 7394 9222
rect 7418 9220 7474 9222
rect 7498 9220 7554 9222
rect 7578 9220 7634 9222
rect 9891 11450 9947 11452
rect 9971 11450 10027 11452
rect 10051 11450 10107 11452
rect 10131 11450 10187 11452
rect 9891 11398 9937 11450
rect 9937 11398 9947 11450
rect 9971 11398 10001 11450
rect 10001 11398 10013 11450
rect 10013 11398 10027 11450
rect 10051 11398 10065 11450
rect 10065 11398 10077 11450
rect 10077 11398 10107 11450
rect 10131 11398 10141 11450
rect 10141 11398 10187 11450
rect 9891 11396 9947 11398
rect 9971 11396 10027 11398
rect 10051 11396 10107 11398
rect 10131 11396 10187 11398
rect 8614 10906 8670 10908
rect 8694 10906 8750 10908
rect 8774 10906 8830 10908
rect 8854 10906 8910 10908
rect 8614 10854 8660 10906
rect 8660 10854 8670 10906
rect 8694 10854 8724 10906
rect 8724 10854 8736 10906
rect 8736 10854 8750 10906
rect 8774 10854 8788 10906
rect 8788 10854 8800 10906
rect 8800 10854 8830 10906
rect 8854 10854 8864 10906
rect 8864 10854 8910 10906
rect 8614 10852 8670 10854
rect 8694 10852 8750 10854
rect 8774 10852 8830 10854
rect 8854 10852 8910 10854
rect 8614 9818 8670 9820
rect 8694 9818 8750 9820
rect 8774 9818 8830 9820
rect 8854 9818 8910 9820
rect 8614 9766 8660 9818
rect 8660 9766 8670 9818
rect 8694 9766 8724 9818
rect 8724 9766 8736 9818
rect 8736 9766 8750 9818
rect 8774 9766 8788 9818
rect 8788 9766 8800 9818
rect 8800 9766 8830 9818
rect 8854 9766 8864 9818
rect 8864 9766 8910 9818
rect 8614 9764 8670 9766
rect 8694 9764 8750 9766
rect 8774 9764 8830 9766
rect 8854 9764 8910 9766
rect 7338 8186 7394 8188
rect 7418 8186 7474 8188
rect 7498 8186 7554 8188
rect 7578 8186 7634 8188
rect 7338 8134 7384 8186
rect 7384 8134 7394 8186
rect 7418 8134 7448 8186
rect 7448 8134 7460 8186
rect 7460 8134 7474 8186
rect 7498 8134 7512 8186
rect 7512 8134 7524 8186
rect 7524 8134 7554 8186
rect 7578 8134 7588 8186
rect 7588 8134 7634 8186
rect 7338 8132 7394 8134
rect 7418 8132 7474 8134
rect 7498 8132 7554 8134
rect 7578 8132 7634 8134
rect 7338 7098 7394 7100
rect 7418 7098 7474 7100
rect 7498 7098 7554 7100
rect 7578 7098 7634 7100
rect 7338 7046 7384 7098
rect 7384 7046 7394 7098
rect 7418 7046 7448 7098
rect 7448 7046 7460 7098
rect 7460 7046 7474 7098
rect 7498 7046 7512 7098
rect 7512 7046 7524 7098
rect 7524 7046 7554 7098
rect 7578 7046 7588 7098
rect 7588 7046 7634 7098
rect 7338 7044 7394 7046
rect 7418 7044 7474 7046
rect 7498 7044 7554 7046
rect 7578 7044 7634 7046
rect 7338 6010 7394 6012
rect 7418 6010 7474 6012
rect 7498 6010 7554 6012
rect 7578 6010 7634 6012
rect 7338 5958 7384 6010
rect 7384 5958 7394 6010
rect 7418 5958 7448 6010
rect 7448 5958 7460 6010
rect 7460 5958 7474 6010
rect 7498 5958 7512 6010
rect 7512 5958 7524 6010
rect 7524 5958 7554 6010
rect 7578 5958 7588 6010
rect 7588 5958 7634 6010
rect 7338 5956 7394 5958
rect 7418 5956 7474 5958
rect 7498 5956 7554 5958
rect 7578 5956 7634 5958
rect 7338 4922 7394 4924
rect 7418 4922 7474 4924
rect 7498 4922 7554 4924
rect 7578 4922 7634 4924
rect 7338 4870 7384 4922
rect 7384 4870 7394 4922
rect 7418 4870 7448 4922
rect 7448 4870 7460 4922
rect 7460 4870 7474 4922
rect 7498 4870 7512 4922
rect 7512 4870 7524 4922
rect 7524 4870 7554 4922
rect 7578 4870 7588 4922
rect 7588 4870 7634 4922
rect 7338 4868 7394 4870
rect 7418 4868 7474 4870
rect 7498 4868 7554 4870
rect 7578 4868 7634 4870
rect 8614 8730 8670 8732
rect 8694 8730 8750 8732
rect 8774 8730 8830 8732
rect 8854 8730 8910 8732
rect 8614 8678 8660 8730
rect 8660 8678 8670 8730
rect 8694 8678 8724 8730
rect 8724 8678 8736 8730
rect 8736 8678 8750 8730
rect 8774 8678 8788 8730
rect 8788 8678 8800 8730
rect 8800 8678 8830 8730
rect 8854 8678 8864 8730
rect 8864 8678 8910 8730
rect 8614 8676 8670 8678
rect 8694 8676 8750 8678
rect 8774 8676 8830 8678
rect 8854 8676 8910 8678
rect 9891 10362 9947 10364
rect 9971 10362 10027 10364
rect 10051 10362 10107 10364
rect 10131 10362 10187 10364
rect 9891 10310 9937 10362
rect 9937 10310 9947 10362
rect 9971 10310 10001 10362
rect 10001 10310 10013 10362
rect 10013 10310 10027 10362
rect 10051 10310 10065 10362
rect 10065 10310 10077 10362
rect 10077 10310 10107 10362
rect 10131 10310 10141 10362
rect 10141 10310 10187 10362
rect 9891 10308 9947 10310
rect 9971 10308 10027 10310
rect 10051 10308 10107 10310
rect 10131 10308 10187 10310
rect 8614 7642 8670 7644
rect 8694 7642 8750 7644
rect 8774 7642 8830 7644
rect 8854 7642 8910 7644
rect 8614 7590 8660 7642
rect 8660 7590 8670 7642
rect 8694 7590 8724 7642
rect 8724 7590 8736 7642
rect 8736 7590 8750 7642
rect 8774 7590 8788 7642
rect 8788 7590 8800 7642
rect 8800 7590 8830 7642
rect 8854 7590 8864 7642
rect 8864 7590 8910 7642
rect 8614 7588 8670 7590
rect 8694 7588 8750 7590
rect 8774 7588 8830 7590
rect 8854 7588 8910 7590
rect 8614 6554 8670 6556
rect 8694 6554 8750 6556
rect 8774 6554 8830 6556
rect 8854 6554 8910 6556
rect 8614 6502 8660 6554
rect 8660 6502 8670 6554
rect 8694 6502 8724 6554
rect 8724 6502 8736 6554
rect 8736 6502 8750 6554
rect 8774 6502 8788 6554
rect 8788 6502 8800 6554
rect 8800 6502 8830 6554
rect 8854 6502 8864 6554
rect 8864 6502 8910 6554
rect 8614 6500 8670 6502
rect 8694 6500 8750 6502
rect 8774 6500 8830 6502
rect 8854 6500 8910 6502
rect 8614 5466 8670 5468
rect 8694 5466 8750 5468
rect 8774 5466 8830 5468
rect 8854 5466 8910 5468
rect 8614 5414 8660 5466
rect 8660 5414 8670 5466
rect 8694 5414 8724 5466
rect 8724 5414 8736 5466
rect 8736 5414 8750 5466
rect 8774 5414 8788 5466
rect 8788 5414 8800 5466
rect 8800 5414 8830 5466
rect 8854 5414 8864 5466
rect 8864 5414 8910 5466
rect 8614 5412 8670 5414
rect 8694 5412 8750 5414
rect 8774 5412 8830 5414
rect 8854 5412 8910 5414
rect 7338 3834 7394 3836
rect 7418 3834 7474 3836
rect 7498 3834 7554 3836
rect 7578 3834 7634 3836
rect 7338 3782 7384 3834
rect 7384 3782 7394 3834
rect 7418 3782 7448 3834
rect 7448 3782 7460 3834
rect 7460 3782 7474 3834
rect 7498 3782 7512 3834
rect 7512 3782 7524 3834
rect 7524 3782 7554 3834
rect 7578 3782 7588 3834
rect 7588 3782 7634 3834
rect 7338 3780 7394 3782
rect 7418 3780 7474 3782
rect 7498 3780 7554 3782
rect 7578 3780 7634 3782
rect 8614 4378 8670 4380
rect 8694 4378 8750 4380
rect 8774 4378 8830 4380
rect 8854 4378 8910 4380
rect 8614 4326 8660 4378
rect 8660 4326 8670 4378
rect 8694 4326 8724 4378
rect 8724 4326 8736 4378
rect 8736 4326 8750 4378
rect 8774 4326 8788 4378
rect 8788 4326 8800 4378
rect 8800 4326 8830 4378
rect 8854 4326 8864 4378
rect 8864 4326 8910 4378
rect 8614 4324 8670 4326
rect 8694 4324 8750 4326
rect 8774 4324 8830 4326
rect 8854 4324 8910 4326
rect 8614 3290 8670 3292
rect 8694 3290 8750 3292
rect 8774 3290 8830 3292
rect 8854 3290 8910 3292
rect 8614 3238 8660 3290
rect 8660 3238 8670 3290
rect 8694 3238 8724 3290
rect 8724 3238 8736 3290
rect 8736 3238 8750 3290
rect 8774 3238 8788 3290
rect 8788 3238 8800 3290
rect 8800 3238 8830 3290
rect 8854 3238 8864 3290
rect 8864 3238 8910 3290
rect 8614 3236 8670 3238
rect 8694 3236 8750 3238
rect 8774 3236 8830 3238
rect 8854 3236 8910 3238
rect 9891 9274 9947 9276
rect 9971 9274 10027 9276
rect 10051 9274 10107 9276
rect 10131 9274 10187 9276
rect 9891 9222 9937 9274
rect 9937 9222 9947 9274
rect 9971 9222 10001 9274
rect 10001 9222 10013 9274
rect 10013 9222 10027 9274
rect 10051 9222 10065 9274
rect 10065 9222 10077 9274
rect 10077 9222 10107 9274
rect 10131 9222 10141 9274
rect 10141 9222 10187 9274
rect 9891 9220 9947 9222
rect 9971 9220 10027 9222
rect 10051 9220 10107 9222
rect 10131 9220 10187 9222
rect 9891 8186 9947 8188
rect 9971 8186 10027 8188
rect 10051 8186 10107 8188
rect 10131 8186 10187 8188
rect 9891 8134 9937 8186
rect 9937 8134 9947 8186
rect 9971 8134 10001 8186
rect 10001 8134 10013 8186
rect 10013 8134 10027 8186
rect 10051 8134 10065 8186
rect 10065 8134 10077 8186
rect 10077 8134 10107 8186
rect 10131 8134 10141 8186
rect 10141 8134 10187 8186
rect 9891 8132 9947 8134
rect 9971 8132 10027 8134
rect 10051 8132 10107 8134
rect 10131 8132 10187 8134
rect 9891 7098 9947 7100
rect 9971 7098 10027 7100
rect 10051 7098 10107 7100
rect 10131 7098 10187 7100
rect 9891 7046 9937 7098
rect 9937 7046 9947 7098
rect 9971 7046 10001 7098
rect 10001 7046 10013 7098
rect 10013 7046 10027 7098
rect 10051 7046 10065 7098
rect 10065 7046 10077 7098
rect 10077 7046 10107 7098
rect 10131 7046 10141 7098
rect 10141 7046 10187 7098
rect 9891 7044 9947 7046
rect 9971 7044 10027 7046
rect 10051 7044 10107 7046
rect 10131 7044 10187 7046
rect 9891 6010 9947 6012
rect 9971 6010 10027 6012
rect 10051 6010 10107 6012
rect 10131 6010 10187 6012
rect 9891 5958 9937 6010
rect 9937 5958 9947 6010
rect 9971 5958 10001 6010
rect 10001 5958 10013 6010
rect 10013 5958 10027 6010
rect 10051 5958 10065 6010
rect 10065 5958 10077 6010
rect 10077 5958 10107 6010
rect 10131 5958 10141 6010
rect 10141 5958 10187 6010
rect 9891 5956 9947 5958
rect 9971 5956 10027 5958
rect 10051 5956 10107 5958
rect 10131 5956 10187 5958
rect 9891 4922 9947 4924
rect 9971 4922 10027 4924
rect 10051 4922 10107 4924
rect 10131 4922 10187 4924
rect 9891 4870 9937 4922
rect 9937 4870 9947 4922
rect 9971 4870 10001 4922
rect 10001 4870 10013 4922
rect 10013 4870 10027 4922
rect 10051 4870 10065 4922
rect 10065 4870 10077 4922
rect 10077 4870 10107 4922
rect 10131 4870 10141 4922
rect 10141 4870 10187 4922
rect 9891 4868 9947 4870
rect 9971 4868 10027 4870
rect 10051 4868 10107 4870
rect 10131 4868 10187 4870
rect 10690 11620 10746 11656
rect 10690 11600 10692 11620
rect 10692 11600 10744 11620
rect 10744 11600 10746 11620
rect 11167 10906 11223 10908
rect 11247 10906 11303 10908
rect 11327 10906 11383 10908
rect 11407 10906 11463 10908
rect 11167 10854 11213 10906
rect 11213 10854 11223 10906
rect 11247 10854 11277 10906
rect 11277 10854 11289 10906
rect 11289 10854 11303 10906
rect 11327 10854 11341 10906
rect 11341 10854 11353 10906
rect 11353 10854 11383 10906
rect 11407 10854 11417 10906
rect 11417 10854 11463 10906
rect 11167 10852 11223 10854
rect 11247 10852 11303 10854
rect 11327 10852 11383 10854
rect 11407 10852 11463 10854
rect 11167 9818 11223 9820
rect 11247 9818 11303 9820
rect 11327 9818 11383 9820
rect 11407 9818 11463 9820
rect 11167 9766 11213 9818
rect 11213 9766 11223 9818
rect 11247 9766 11277 9818
rect 11277 9766 11289 9818
rect 11289 9766 11303 9818
rect 11327 9766 11341 9818
rect 11341 9766 11353 9818
rect 11353 9766 11383 9818
rect 11407 9766 11417 9818
rect 11417 9766 11463 9818
rect 11167 9764 11223 9766
rect 11247 9764 11303 9766
rect 11327 9764 11383 9766
rect 11407 9764 11463 9766
rect 11167 8730 11223 8732
rect 11247 8730 11303 8732
rect 11327 8730 11383 8732
rect 11407 8730 11463 8732
rect 11167 8678 11213 8730
rect 11213 8678 11223 8730
rect 11247 8678 11277 8730
rect 11277 8678 11289 8730
rect 11289 8678 11303 8730
rect 11327 8678 11341 8730
rect 11341 8678 11353 8730
rect 11353 8678 11383 8730
rect 11407 8678 11417 8730
rect 11417 8678 11463 8730
rect 11167 8676 11223 8678
rect 11247 8676 11303 8678
rect 11327 8676 11383 8678
rect 11407 8676 11463 8678
rect 11167 7642 11223 7644
rect 11247 7642 11303 7644
rect 11327 7642 11383 7644
rect 11407 7642 11463 7644
rect 11167 7590 11213 7642
rect 11213 7590 11223 7642
rect 11247 7590 11277 7642
rect 11277 7590 11289 7642
rect 11289 7590 11303 7642
rect 11327 7590 11341 7642
rect 11341 7590 11353 7642
rect 11353 7590 11383 7642
rect 11407 7590 11417 7642
rect 11417 7590 11463 7642
rect 11167 7588 11223 7590
rect 11247 7588 11303 7590
rect 11327 7588 11383 7590
rect 11407 7588 11463 7590
rect 11167 6554 11223 6556
rect 11247 6554 11303 6556
rect 11327 6554 11383 6556
rect 11407 6554 11463 6556
rect 11167 6502 11213 6554
rect 11213 6502 11223 6554
rect 11247 6502 11277 6554
rect 11277 6502 11289 6554
rect 11289 6502 11303 6554
rect 11327 6502 11341 6554
rect 11341 6502 11353 6554
rect 11353 6502 11383 6554
rect 11407 6502 11417 6554
rect 11417 6502 11463 6554
rect 11167 6500 11223 6502
rect 11247 6500 11303 6502
rect 11327 6500 11383 6502
rect 11407 6500 11463 6502
rect 11167 5466 11223 5468
rect 11247 5466 11303 5468
rect 11327 5466 11383 5468
rect 11407 5466 11463 5468
rect 11167 5414 11213 5466
rect 11213 5414 11223 5466
rect 11247 5414 11277 5466
rect 11277 5414 11289 5466
rect 11289 5414 11303 5466
rect 11327 5414 11341 5466
rect 11341 5414 11353 5466
rect 11353 5414 11383 5466
rect 11407 5414 11417 5466
rect 11417 5414 11463 5466
rect 11167 5412 11223 5414
rect 11247 5412 11303 5414
rect 11327 5412 11383 5414
rect 11407 5412 11463 5414
rect 10782 5208 10838 5264
rect 11167 4378 11223 4380
rect 11247 4378 11303 4380
rect 11327 4378 11383 4380
rect 11407 4378 11463 4380
rect 11167 4326 11213 4378
rect 11213 4326 11223 4378
rect 11247 4326 11277 4378
rect 11277 4326 11289 4378
rect 11289 4326 11303 4378
rect 11327 4326 11341 4378
rect 11341 4326 11353 4378
rect 11353 4326 11383 4378
rect 11407 4326 11417 4378
rect 11417 4326 11463 4378
rect 11167 4324 11223 4326
rect 11247 4324 11303 4326
rect 11327 4324 11383 4326
rect 11407 4324 11463 4326
rect 9891 3834 9947 3836
rect 9971 3834 10027 3836
rect 10051 3834 10107 3836
rect 10131 3834 10187 3836
rect 9891 3782 9937 3834
rect 9937 3782 9947 3834
rect 9971 3782 10001 3834
rect 10001 3782 10013 3834
rect 10013 3782 10027 3834
rect 10051 3782 10065 3834
rect 10065 3782 10077 3834
rect 10077 3782 10107 3834
rect 10131 3782 10141 3834
rect 10141 3782 10187 3834
rect 9891 3780 9947 3782
rect 9971 3780 10027 3782
rect 10051 3780 10107 3782
rect 10131 3780 10187 3782
rect 11167 3290 11223 3292
rect 11247 3290 11303 3292
rect 11327 3290 11383 3292
rect 11407 3290 11463 3292
rect 11167 3238 11213 3290
rect 11213 3238 11223 3290
rect 11247 3238 11277 3290
rect 11277 3238 11289 3290
rect 11289 3238 11303 3290
rect 11327 3238 11341 3290
rect 11341 3238 11353 3290
rect 11353 3238 11383 3290
rect 11407 3238 11417 3290
rect 11417 3238 11463 3290
rect 11167 3236 11223 3238
rect 11247 3236 11303 3238
rect 11327 3236 11383 3238
rect 11407 3236 11463 3238
rect 7338 2746 7394 2748
rect 7418 2746 7474 2748
rect 7498 2746 7554 2748
rect 7578 2746 7634 2748
rect 7338 2694 7384 2746
rect 7384 2694 7394 2746
rect 7418 2694 7448 2746
rect 7448 2694 7460 2746
rect 7460 2694 7474 2746
rect 7498 2694 7512 2746
rect 7512 2694 7524 2746
rect 7524 2694 7554 2746
rect 7578 2694 7588 2746
rect 7588 2694 7634 2746
rect 7338 2692 7394 2694
rect 7418 2692 7474 2694
rect 7498 2692 7554 2694
rect 7578 2692 7634 2694
rect 9891 2746 9947 2748
rect 9971 2746 10027 2748
rect 10051 2746 10107 2748
rect 10131 2746 10187 2748
rect 9891 2694 9937 2746
rect 9937 2694 9947 2746
rect 9971 2694 10001 2746
rect 10001 2694 10013 2746
rect 10013 2694 10027 2746
rect 10051 2694 10065 2746
rect 10065 2694 10077 2746
rect 10077 2694 10107 2746
rect 10131 2694 10141 2746
rect 10141 2694 10187 2746
rect 9891 2692 9947 2694
rect 9971 2692 10027 2694
rect 10051 2692 10107 2694
rect 10131 2692 10187 2694
rect 3508 2202 3564 2204
rect 3588 2202 3644 2204
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3508 2150 3554 2202
rect 3554 2150 3564 2202
rect 3588 2150 3618 2202
rect 3618 2150 3630 2202
rect 3630 2150 3644 2202
rect 3668 2150 3682 2202
rect 3682 2150 3694 2202
rect 3694 2150 3724 2202
rect 3748 2150 3758 2202
rect 3758 2150 3804 2202
rect 3508 2148 3564 2150
rect 3588 2148 3644 2150
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 6061 2202 6117 2204
rect 6141 2202 6197 2204
rect 6221 2202 6277 2204
rect 6301 2202 6357 2204
rect 6061 2150 6107 2202
rect 6107 2150 6117 2202
rect 6141 2150 6171 2202
rect 6171 2150 6183 2202
rect 6183 2150 6197 2202
rect 6221 2150 6235 2202
rect 6235 2150 6247 2202
rect 6247 2150 6277 2202
rect 6301 2150 6311 2202
rect 6311 2150 6357 2202
rect 6061 2148 6117 2150
rect 6141 2148 6197 2150
rect 6221 2148 6277 2150
rect 6301 2148 6357 2150
rect 8614 2202 8670 2204
rect 8694 2202 8750 2204
rect 8774 2202 8830 2204
rect 8854 2202 8910 2204
rect 8614 2150 8660 2202
rect 8660 2150 8670 2202
rect 8694 2150 8724 2202
rect 8724 2150 8736 2202
rect 8736 2150 8750 2202
rect 8774 2150 8788 2202
rect 8788 2150 8800 2202
rect 8800 2150 8830 2202
rect 8854 2150 8864 2202
rect 8864 2150 8910 2202
rect 8614 2148 8670 2150
rect 8694 2148 8750 2150
rect 8774 2148 8830 2150
rect 8854 2148 8910 2150
rect 11167 2202 11223 2204
rect 11247 2202 11303 2204
rect 11327 2202 11383 2204
rect 11407 2202 11463 2204
rect 11167 2150 11213 2202
rect 11213 2150 11223 2202
rect 11247 2150 11277 2202
rect 11277 2150 11289 2202
rect 11289 2150 11303 2202
rect 11327 2150 11341 2202
rect 11341 2150 11353 2202
rect 11353 2150 11383 2202
rect 11407 2150 11417 2202
rect 11417 2150 11463 2202
rect 11167 2148 11223 2150
rect 11247 2148 11303 2150
rect 11327 2148 11383 2150
rect 11407 2148 11463 2150
<< metal3 >>
rect 0 12338 800 12368
rect 1669 12338 1735 12341
rect 0 12336 1735 12338
rect 0 12280 1674 12336
rect 1730 12280 1735 12336
rect 0 12278 1735 12280
rect 0 12248 800 12278
rect 1669 12275 1735 12278
rect 3498 12000 3814 12001
rect 3498 11936 3504 12000
rect 3568 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3814 12000
rect 3498 11935 3814 11936
rect 6051 12000 6367 12001
rect 6051 11936 6057 12000
rect 6121 11936 6137 12000
rect 6201 11936 6217 12000
rect 6281 11936 6297 12000
rect 6361 11936 6367 12000
rect 6051 11935 6367 11936
rect 8604 12000 8920 12001
rect 8604 11936 8610 12000
rect 8674 11936 8690 12000
rect 8754 11936 8770 12000
rect 8834 11936 8850 12000
rect 8914 11936 8920 12000
rect 8604 11935 8920 11936
rect 11157 12000 11473 12001
rect 11157 11936 11163 12000
rect 11227 11936 11243 12000
rect 11307 11936 11323 12000
rect 11387 11936 11403 12000
rect 11467 11936 11473 12000
rect 11157 11935 11473 11936
rect 10685 11658 10751 11661
rect 11708 11658 12508 11688
rect 10685 11656 12508 11658
rect 10685 11600 10690 11656
rect 10746 11600 12508 11656
rect 10685 11598 12508 11600
rect 10685 11595 10751 11598
rect 11708 11568 12508 11598
rect 2222 11456 2538 11457
rect 2222 11392 2228 11456
rect 2292 11392 2308 11456
rect 2372 11392 2388 11456
rect 2452 11392 2468 11456
rect 2532 11392 2538 11456
rect 2222 11391 2538 11392
rect 4775 11456 5091 11457
rect 4775 11392 4781 11456
rect 4845 11392 4861 11456
rect 4925 11392 4941 11456
rect 5005 11392 5021 11456
rect 5085 11392 5091 11456
rect 4775 11391 5091 11392
rect 7328 11456 7644 11457
rect 7328 11392 7334 11456
rect 7398 11392 7414 11456
rect 7478 11392 7494 11456
rect 7558 11392 7574 11456
rect 7638 11392 7644 11456
rect 7328 11391 7644 11392
rect 9881 11456 10197 11457
rect 9881 11392 9887 11456
rect 9951 11392 9967 11456
rect 10031 11392 10047 11456
rect 10111 11392 10127 11456
rect 10191 11392 10197 11456
rect 9881 11391 10197 11392
rect 3498 10912 3814 10913
rect 3498 10848 3504 10912
rect 3568 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3814 10912
rect 3498 10847 3814 10848
rect 6051 10912 6367 10913
rect 6051 10848 6057 10912
rect 6121 10848 6137 10912
rect 6201 10848 6217 10912
rect 6281 10848 6297 10912
rect 6361 10848 6367 10912
rect 6051 10847 6367 10848
rect 8604 10912 8920 10913
rect 8604 10848 8610 10912
rect 8674 10848 8690 10912
rect 8754 10848 8770 10912
rect 8834 10848 8850 10912
rect 8914 10848 8920 10912
rect 8604 10847 8920 10848
rect 11157 10912 11473 10913
rect 11157 10848 11163 10912
rect 11227 10848 11243 10912
rect 11307 10848 11323 10912
rect 11387 10848 11403 10912
rect 11467 10848 11473 10912
rect 11157 10847 11473 10848
rect 2222 10368 2538 10369
rect 2222 10304 2228 10368
rect 2292 10304 2308 10368
rect 2372 10304 2388 10368
rect 2452 10304 2468 10368
rect 2532 10304 2538 10368
rect 2222 10303 2538 10304
rect 4775 10368 5091 10369
rect 4775 10304 4781 10368
rect 4845 10304 4861 10368
rect 4925 10304 4941 10368
rect 5005 10304 5021 10368
rect 5085 10304 5091 10368
rect 4775 10303 5091 10304
rect 7328 10368 7644 10369
rect 7328 10304 7334 10368
rect 7398 10304 7414 10368
rect 7478 10304 7494 10368
rect 7558 10304 7574 10368
rect 7638 10304 7644 10368
rect 7328 10303 7644 10304
rect 9881 10368 10197 10369
rect 9881 10304 9887 10368
rect 9951 10304 9967 10368
rect 10031 10304 10047 10368
rect 10111 10304 10127 10368
rect 10191 10304 10197 10368
rect 9881 10303 10197 10304
rect 3498 9824 3814 9825
rect 3498 9760 3504 9824
rect 3568 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3814 9824
rect 3498 9759 3814 9760
rect 6051 9824 6367 9825
rect 6051 9760 6057 9824
rect 6121 9760 6137 9824
rect 6201 9760 6217 9824
rect 6281 9760 6297 9824
rect 6361 9760 6367 9824
rect 6051 9759 6367 9760
rect 8604 9824 8920 9825
rect 8604 9760 8610 9824
rect 8674 9760 8690 9824
rect 8754 9760 8770 9824
rect 8834 9760 8850 9824
rect 8914 9760 8920 9824
rect 8604 9759 8920 9760
rect 11157 9824 11473 9825
rect 11157 9760 11163 9824
rect 11227 9760 11243 9824
rect 11307 9760 11323 9824
rect 11387 9760 11403 9824
rect 11467 9760 11473 9824
rect 11157 9759 11473 9760
rect 2222 9280 2538 9281
rect 2222 9216 2228 9280
rect 2292 9216 2308 9280
rect 2372 9216 2388 9280
rect 2452 9216 2468 9280
rect 2532 9216 2538 9280
rect 2222 9215 2538 9216
rect 4775 9280 5091 9281
rect 4775 9216 4781 9280
rect 4845 9216 4861 9280
rect 4925 9216 4941 9280
rect 5005 9216 5021 9280
rect 5085 9216 5091 9280
rect 4775 9215 5091 9216
rect 7328 9280 7644 9281
rect 7328 9216 7334 9280
rect 7398 9216 7414 9280
rect 7478 9216 7494 9280
rect 7558 9216 7574 9280
rect 7638 9216 7644 9280
rect 7328 9215 7644 9216
rect 9881 9280 10197 9281
rect 9881 9216 9887 9280
rect 9951 9216 9967 9280
rect 10031 9216 10047 9280
rect 10111 9216 10127 9280
rect 10191 9216 10197 9280
rect 9881 9215 10197 9216
rect 3498 8736 3814 8737
rect 3498 8672 3504 8736
rect 3568 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3814 8736
rect 3498 8671 3814 8672
rect 6051 8736 6367 8737
rect 6051 8672 6057 8736
rect 6121 8672 6137 8736
rect 6201 8672 6217 8736
rect 6281 8672 6297 8736
rect 6361 8672 6367 8736
rect 6051 8671 6367 8672
rect 8604 8736 8920 8737
rect 8604 8672 8610 8736
rect 8674 8672 8690 8736
rect 8754 8672 8770 8736
rect 8834 8672 8850 8736
rect 8914 8672 8920 8736
rect 8604 8671 8920 8672
rect 11157 8736 11473 8737
rect 11157 8672 11163 8736
rect 11227 8672 11243 8736
rect 11307 8672 11323 8736
rect 11387 8672 11403 8736
rect 11467 8672 11473 8736
rect 11157 8671 11473 8672
rect 2222 8192 2538 8193
rect 2222 8128 2228 8192
rect 2292 8128 2308 8192
rect 2372 8128 2388 8192
rect 2452 8128 2468 8192
rect 2532 8128 2538 8192
rect 2222 8127 2538 8128
rect 4775 8192 5091 8193
rect 4775 8128 4781 8192
rect 4845 8128 4861 8192
rect 4925 8128 4941 8192
rect 5005 8128 5021 8192
rect 5085 8128 5091 8192
rect 4775 8127 5091 8128
rect 7328 8192 7644 8193
rect 7328 8128 7334 8192
rect 7398 8128 7414 8192
rect 7478 8128 7494 8192
rect 7558 8128 7574 8192
rect 7638 8128 7644 8192
rect 7328 8127 7644 8128
rect 9881 8192 10197 8193
rect 9881 8128 9887 8192
rect 9951 8128 9967 8192
rect 10031 8128 10047 8192
rect 10111 8128 10127 8192
rect 10191 8128 10197 8192
rect 9881 8127 10197 8128
rect 3498 7648 3814 7649
rect 3498 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3814 7648
rect 3498 7583 3814 7584
rect 6051 7648 6367 7649
rect 6051 7584 6057 7648
rect 6121 7584 6137 7648
rect 6201 7584 6217 7648
rect 6281 7584 6297 7648
rect 6361 7584 6367 7648
rect 6051 7583 6367 7584
rect 8604 7648 8920 7649
rect 8604 7584 8610 7648
rect 8674 7584 8690 7648
rect 8754 7584 8770 7648
rect 8834 7584 8850 7648
rect 8914 7584 8920 7648
rect 8604 7583 8920 7584
rect 11157 7648 11473 7649
rect 11157 7584 11163 7648
rect 11227 7584 11243 7648
rect 11307 7584 11323 7648
rect 11387 7584 11403 7648
rect 11467 7584 11473 7648
rect 11157 7583 11473 7584
rect 2222 7104 2538 7105
rect 2222 7040 2228 7104
rect 2292 7040 2308 7104
rect 2372 7040 2388 7104
rect 2452 7040 2468 7104
rect 2532 7040 2538 7104
rect 2222 7039 2538 7040
rect 4775 7104 5091 7105
rect 4775 7040 4781 7104
rect 4845 7040 4861 7104
rect 4925 7040 4941 7104
rect 5005 7040 5021 7104
rect 5085 7040 5091 7104
rect 4775 7039 5091 7040
rect 7328 7104 7644 7105
rect 7328 7040 7334 7104
rect 7398 7040 7414 7104
rect 7478 7040 7494 7104
rect 7558 7040 7574 7104
rect 7638 7040 7644 7104
rect 7328 7039 7644 7040
rect 9881 7104 10197 7105
rect 9881 7040 9887 7104
rect 9951 7040 9967 7104
rect 10031 7040 10047 7104
rect 10111 7040 10127 7104
rect 10191 7040 10197 7104
rect 9881 7039 10197 7040
rect 3498 6560 3814 6561
rect 3498 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3814 6560
rect 3498 6495 3814 6496
rect 6051 6560 6367 6561
rect 6051 6496 6057 6560
rect 6121 6496 6137 6560
rect 6201 6496 6217 6560
rect 6281 6496 6297 6560
rect 6361 6496 6367 6560
rect 6051 6495 6367 6496
rect 8604 6560 8920 6561
rect 8604 6496 8610 6560
rect 8674 6496 8690 6560
rect 8754 6496 8770 6560
rect 8834 6496 8850 6560
rect 8914 6496 8920 6560
rect 8604 6495 8920 6496
rect 11157 6560 11473 6561
rect 11157 6496 11163 6560
rect 11227 6496 11243 6560
rect 11307 6496 11323 6560
rect 11387 6496 11403 6560
rect 11467 6496 11473 6560
rect 11157 6495 11473 6496
rect 0 6128 800 6248
rect 2222 6016 2538 6017
rect 2222 5952 2228 6016
rect 2292 5952 2308 6016
rect 2372 5952 2388 6016
rect 2452 5952 2468 6016
rect 2532 5952 2538 6016
rect 2222 5951 2538 5952
rect 4775 6016 5091 6017
rect 4775 5952 4781 6016
rect 4845 5952 4861 6016
rect 4925 5952 4941 6016
rect 5005 5952 5021 6016
rect 5085 5952 5091 6016
rect 4775 5951 5091 5952
rect 7328 6016 7644 6017
rect 7328 5952 7334 6016
rect 7398 5952 7414 6016
rect 7478 5952 7494 6016
rect 7558 5952 7574 6016
rect 7638 5952 7644 6016
rect 7328 5951 7644 5952
rect 9881 6016 10197 6017
rect 9881 5952 9887 6016
rect 9951 5952 9967 6016
rect 10031 5952 10047 6016
rect 10111 5952 10127 6016
rect 10191 5952 10197 6016
rect 9881 5951 10197 5952
rect 11708 5538 12508 5568
rect 3498 5472 3814 5473
rect 3498 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3814 5472
rect 3498 5407 3814 5408
rect 6051 5472 6367 5473
rect 6051 5408 6057 5472
rect 6121 5408 6137 5472
rect 6201 5408 6217 5472
rect 6281 5408 6297 5472
rect 6361 5408 6367 5472
rect 6051 5407 6367 5408
rect 8604 5472 8920 5473
rect 8604 5408 8610 5472
rect 8674 5408 8690 5472
rect 8754 5408 8770 5472
rect 8834 5408 8850 5472
rect 8914 5408 8920 5472
rect 8604 5407 8920 5408
rect 11157 5472 11473 5473
rect 11157 5408 11163 5472
rect 11227 5408 11243 5472
rect 11307 5408 11323 5472
rect 11387 5408 11403 5472
rect 11467 5408 11473 5472
rect 11157 5407 11473 5408
rect 11654 5448 12508 5538
rect 10777 5266 10843 5269
rect 11654 5266 11714 5448
rect 10777 5264 11714 5266
rect 10777 5208 10782 5264
rect 10838 5208 11714 5264
rect 10777 5206 11714 5208
rect 10777 5203 10843 5206
rect 2222 4928 2538 4929
rect 2222 4864 2228 4928
rect 2292 4864 2308 4928
rect 2372 4864 2388 4928
rect 2452 4864 2468 4928
rect 2532 4864 2538 4928
rect 2222 4863 2538 4864
rect 4775 4928 5091 4929
rect 4775 4864 4781 4928
rect 4845 4864 4861 4928
rect 4925 4864 4941 4928
rect 5005 4864 5021 4928
rect 5085 4864 5091 4928
rect 4775 4863 5091 4864
rect 7328 4928 7644 4929
rect 7328 4864 7334 4928
rect 7398 4864 7414 4928
rect 7478 4864 7494 4928
rect 7558 4864 7574 4928
rect 7638 4864 7644 4928
rect 7328 4863 7644 4864
rect 9881 4928 10197 4929
rect 9881 4864 9887 4928
rect 9951 4864 9967 4928
rect 10031 4864 10047 4928
rect 10111 4864 10127 4928
rect 10191 4864 10197 4928
rect 9881 4863 10197 4864
rect 3498 4384 3814 4385
rect 3498 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3814 4384
rect 3498 4319 3814 4320
rect 6051 4384 6367 4385
rect 6051 4320 6057 4384
rect 6121 4320 6137 4384
rect 6201 4320 6217 4384
rect 6281 4320 6297 4384
rect 6361 4320 6367 4384
rect 6051 4319 6367 4320
rect 8604 4384 8920 4385
rect 8604 4320 8610 4384
rect 8674 4320 8690 4384
rect 8754 4320 8770 4384
rect 8834 4320 8850 4384
rect 8914 4320 8920 4384
rect 8604 4319 8920 4320
rect 11157 4384 11473 4385
rect 11157 4320 11163 4384
rect 11227 4320 11243 4384
rect 11307 4320 11323 4384
rect 11387 4320 11403 4384
rect 11467 4320 11473 4384
rect 11157 4319 11473 4320
rect 2222 3840 2538 3841
rect 2222 3776 2228 3840
rect 2292 3776 2308 3840
rect 2372 3776 2388 3840
rect 2452 3776 2468 3840
rect 2532 3776 2538 3840
rect 2222 3775 2538 3776
rect 4775 3840 5091 3841
rect 4775 3776 4781 3840
rect 4845 3776 4861 3840
rect 4925 3776 4941 3840
rect 5005 3776 5021 3840
rect 5085 3776 5091 3840
rect 4775 3775 5091 3776
rect 7328 3840 7644 3841
rect 7328 3776 7334 3840
rect 7398 3776 7414 3840
rect 7478 3776 7494 3840
rect 7558 3776 7574 3840
rect 7638 3776 7644 3840
rect 7328 3775 7644 3776
rect 9881 3840 10197 3841
rect 9881 3776 9887 3840
rect 9951 3776 9967 3840
rect 10031 3776 10047 3840
rect 10111 3776 10127 3840
rect 10191 3776 10197 3840
rect 9881 3775 10197 3776
rect 3498 3296 3814 3297
rect 3498 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3814 3296
rect 3498 3231 3814 3232
rect 6051 3296 6367 3297
rect 6051 3232 6057 3296
rect 6121 3232 6137 3296
rect 6201 3232 6217 3296
rect 6281 3232 6297 3296
rect 6361 3232 6367 3296
rect 6051 3231 6367 3232
rect 8604 3296 8920 3297
rect 8604 3232 8610 3296
rect 8674 3232 8690 3296
rect 8754 3232 8770 3296
rect 8834 3232 8850 3296
rect 8914 3232 8920 3296
rect 8604 3231 8920 3232
rect 11157 3296 11473 3297
rect 11157 3232 11163 3296
rect 11227 3232 11243 3296
rect 11307 3232 11323 3296
rect 11387 3232 11403 3296
rect 11467 3232 11473 3296
rect 11157 3231 11473 3232
rect 2222 2752 2538 2753
rect 2222 2688 2228 2752
rect 2292 2688 2308 2752
rect 2372 2688 2388 2752
rect 2452 2688 2468 2752
rect 2532 2688 2538 2752
rect 2222 2687 2538 2688
rect 4775 2752 5091 2753
rect 4775 2688 4781 2752
rect 4845 2688 4861 2752
rect 4925 2688 4941 2752
rect 5005 2688 5021 2752
rect 5085 2688 5091 2752
rect 4775 2687 5091 2688
rect 7328 2752 7644 2753
rect 7328 2688 7334 2752
rect 7398 2688 7414 2752
rect 7478 2688 7494 2752
rect 7558 2688 7574 2752
rect 7638 2688 7644 2752
rect 7328 2687 7644 2688
rect 9881 2752 10197 2753
rect 9881 2688 9887 2752
rect 9951 2688 9967 2752
rect 10031 2688 10047 2752
rect 10111 2688 10127 2752
rect 10191 2688 10197 2752
rect 9881 2687 10197 2688
rect 3498 2208 3814 2209
rect 3498 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3814 2208
rect 3498 2143 3814 2144
rect 6051 2208 6367 2209
rect 6051 2144 6057 2208
rect 6121 2144 6137 2208
rect 6201 2144 6217 2208
rect 6281 2144 6297 2208
rect 6361 2144 6367 2208
rect 6051 2143 6367 2144
rect 8604 2208 8920 2209
rect 8604 2144 8610 2208
rect 8674 2144 8690 2208
rect 8754 2144 8770 2208
rect 8834 2144 8850 2208
rect 8914 2144 8920 2208
rect 8604 2143 8920 2144
rect 11157 2208 11473 2209
rect 11157 2144 11163 2208
rect 11227 2144 11243 2208
rect 11307 2144 11323 2208
rect 11387 2144 11403 2208
rect 11467 2144 11473 2208
rect 11157 2143 11473 2144
<< via3 >>
rect 3504 11996 3568 12000
rect 3504 11940 3508 11996
rect 3508 11940 3564 11996
rect 3564 11940 3568 11996
rect 3504 11936 3568 11940
rect 3584 11996 3648 12000
rect 3584 11940 3588 11996
rect 3588 11940 3644 11996
rect 3644 11940 3648 11996
rect 3584 11936 3648 11940
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 6057 11996 6121 12000
rect 6057 11940 6061 11996
rect 6061 11940 6117 11996
rect 6117 11940 6121 11996
rect 6057 11936 6121 11940
rect 6137 11996 6201 12000
rect 6137 11940 6141 11996
rect 6141 11940 6197 11996
rect 6197 11940 6201 11996
rect 6137 11936 6201 11940
rect 6217 11996 6281 12000
rect 6217 11940 6221 11996
rect 6221 11940 6277 11996
rect 6277 11940 6281 11996
rect 6217 11936 6281 11940
rect 6297 11996 6361 12000
rect 6297 11940 6301 11996
rect 6301 11940 6357 11996
rect 6357 11940 6361 11996
rect 6297 11936 6361 11940
rect 8610 11996 8674 12000
rect 8610 11940 8614 11996
rect 8614 11940 8670 11996
rect 8670 11940 8674 11996
rect 8610 11936 8674 11940
rect 8690 11996 8754 12000
rect 8690 11940 8694 11996
rect 8694 11940 8750 11996
rect 8750 11940 8754 11996
rect 8690 11936 8754 11940
rect 8770 11996 8834 12000
rect 8770 11940 8774 11996
rect 8774 11940 8830 11996
rect 8830 11940 8834 11996
rect 8770 11936 8834 11940
rect 8850 11996 8914 12000
rect 8850 11940 8854 11996
rect 8854 11940 8910 11996
rect 8910 11940 8914 11996
rect 8850 11936 8914 11940
rect 11163 11996 11227 12000
rect 11163 11940 11167 11996
rect 11167 11940 11223 11996
rect 11223 11940 11227 11996
rect 11163 11936 11227 11940
rect 11243 11996 11307 12000
rect 11243 11940 11247 11996
rect 11247 11940 11303 11996
rect 11303 11940 11307 11996
rect 11243 11936 11307 11940
rect 11323 11996 11387 12000
rect 11323 11940 11327 11996
rect 11327 11940 11383 11996
rect 11383 11940 11387 11996
rect 11323 11936 11387 11940
rect 11403 11996 11467 12000
rect 11403 11940 11407 11996
rect 11407 11940 11463 11996
rect 11463 11940 11467 11996
rect 11403 11936 11467 11940
rect 2228 11452 2292 11456
rect 2228 11396 2232 11452
rect 2232 11396 2288 11452
rect 2288 11396 2292 11452
rect 2228 11392 2292 11396
rect 2308 11452 2372 11456
rect 2308 11396 2312 11452
rect 2312 11396 2368 11452
rect 2368 11396 2372 11452
rect 2308 11392 2372 11396
rect 2388 11452 2452 11456
rect 2388 11396 2392 11452
rect 2392 11396 2448 11452
rect 2448 11396 2452 11452
rect 2388 11392 2452 11396
rect 2468 11452 2532 11456
rect 2468 11396 2472 11452
rect 2472 11396 2528 11452
rect 2528 11396 2532 11452
rect 2468 11392 2532 11396
rect 4781 11452 4845 11456
rect 4781 11396 4785 11452
rect 4785 11396 4841 11452
rect 4841 11396 4845 11452
rect 4781 11392 4845 11396
rect 4861 11452 4925 11456
rect 4861 11396 4865 11452
rect 4865 11396 4921 11452
rect 4921 11396 4925 11452
rect 4861 11392 4925 11396
rect 4941 11452 5005 11456
rect 4941 11396 4945 11452
rect 4945 11396 5001 11452
rect 5001 11396 5005 11452
rect 4941 11392 5005 11396
rect 5021 11452 5085 11456
rect 5021 11396 5025 11452
rect 5025 11396 5081 11452
rect 5081 11396 5085 11452
rect 5021 11392 5085 11396
rect 7334 11452 7398 11456
rect 7334 11396 7338 11452
rect 7338 11396 7394 11452
rect 7394 11396 7398 11452
rect 7334 11392 7398 11396
rect 7414 11452 7478 11456
rect 7414 11396 7418 11452
rect 7418 11396 7474 11452
rect 7474 11396 7478 11452
rect 7414 11392 7478 11396
rect 7494 11452 7558 11456
rect 7494 11396 7498 11452
rect 7498 11396 7554 11452
rect 7554 11396 7558 11452
rect 7494 11392 7558 11396
rect 7574 11452 7638 11456
rect 7574 11396 7578 11452
rect 7578 11396 7634 11452
rect 7634 11396 7638 11452
rect 7574 11392 7638 11396
rect 9887 11452 9951 11456
rect 9887 11396 9891 11452
rect 9891 11396 9947 11452
rect 9947 11396 9951 11452
rect 9887 11392 9951 11396
rect 9967 11452 10031 11456
rect 9967 11396 9971 11452
rect 9971 11396 10027 11452
rect 10027 11396 10031 11452
rect 9967 11392 10031 11396
rect 10047 11452 10111 11456
rect 10047 11396 10051 11452
rect 10051 11396 10107 11452
rect 10107 11396 10111 11452
rect 10047 11392 10111 11396
rect 10127 11452 10191 11456
rect 10127 11396 10131 11452
rect 10131 11396 10187 11452
rect 10187 11396 10191 11452
rect 10127 11392 10191 11396
rect 3504 10908 3568 10912
rect 3504 10852 3508 10908
rect 3508 10852 3564 10908
rect 3564 10852 3568 10908
rect 3504 10848 3568 10852
rect 3584 10908 3648 10912
rect 3584 10852 3588 10908
rect 3588 10852 3644 10908
rect 3644 10852 3648 10908
rect 3584 10848 3648 10852
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 6057 10908 6121 10912
rect 6057 10852 6061 10908
rect 6061 10852 6117 10908
rect 6117 10852 6121 10908
rect 6057 10848 6121 10852
rect 6137 10908 6201 10912
rect 6137 10852 6141 10908
rect 6141 10852 6197 10908
rect 6197 10852 6201 10908
rect 6137 10848 6201 10852
rect 6217 10908 6281 10912
rect 6217 10852 6221 10908
rect 6221 10852 6277 10908
rect 6277 10852 6281 10908
rect 6217 10848 6281 10852
rect 6297 10908 6361 10912
rect 6297 10852 6301 10908
rect 6301 10852 6357 10908
rect 6357 10852 6361 10908
rect 6297 10848 6361 10852
rect 8610 10908 8674 10912
rect 8610 10852 8614 10908
rect 8614 10852 8670 10908
rect 8670 10852 8674 10908
rect 8610 10848 8674 10852
rect 8690 10908 8754 10912
rect 8690 10852 8694 10908
rect 8694 10852 8750 10908
rect 8750 10852 8754 10908
rect 8690 10848 8754 10852
rect 8770 10908 8834 10912
rect 8770 10852 8774 10908
rect 8774 10852 8830 10908
rect 8830 10852 8834 10908
rect 8770 10848 8834 10852
rect 8850 10908 8914 10912
rect 8850 10852 8854 10908
rect 8854 10852 8910 10908
rect 8910 10852 8914 10908
rect 8850 10848 8914 10852
rect 11163 10908 11227 10912
rect 11163 10852 11167 10908
rect 11167 10852 11223 10908
rect 11223 10852 11227 10908
rect 11163 10848 11227 10852
rect 11243 10908 11307 10912
rect 11243 10852 11247 10908
rect 11247 10852 11303 10908
rect 11303 10852 11307 10908
rect 11243 10848 11307 10852
rect 11323 10908 11387 10912
rect 11323 10852 11327 10908
rect 11327 10852 11383 10908
rect 11383 10852 11387 10908
rect 11323 10848 11387 10852
rect 11403 10908 11467 10912
rect 11403 10852 11407 10908
rect 11407 10852 11463 10908
rect 11463 10852 11467 10908
rect 11403 10848 11467 10852
rect 2228 10364 2292 10368
rect 2228 10308 2232 10364
rect 2232 10308 2288 10364
rect 2288 10308 2292 10364
rect 2228 10304 2292 10308
rect 2308 10364 2372 10368
rect 2308 10308 2312 10364
rect 2312 10308 2368 10364
rect 2368 10308 2372 10364
rect 2308 10304 2372 10308
rect 2388 10364 2452 10368
rect 2388 10308 2392 10364
rect 2392 10308 2448 10364
rect 2448 10308 2452 10364
rect 2388 10304 2452 10308
rect 2468 10364 2532 10368
rect 2468 10308 2472 10364
rect 2472 10308 2528 10364
rect 2528 10308 2532 10364
rect 2468 10304 2532 10308
rect 4781 10364 4845 10368
rect 4781 10308 4785 10364
rect 4785 10308 4841 10364
rect 4841 10308 4845 10364
rect 4781 10304 4845 10308
rect 4861 10364 4925 10368
rect 4861 10308 4865 10364
rect 4865 10308 4921 10364
rect 4921 10308 4925 10364
rect 4861 10304 4925 10308
rect 4941 10364 5005 10368
rect 4941 10308 4945 10364
rect 4945 10308 5001 10364
rect 5001 10308 5005 10364
rect 4941 10304 5005 10308
rect 5021 10364 5085 10368
rect 5021 10308 5025 10364
rect 5025 10308 5081 10364
rect 5081 10308 5085 10364
rect 5021 10304 5085 10308
rect 7334 10364 7398 10368
rect 7334 10308 7338 10364
rect 7338 10308 7394 10364
rect 7394 10308 7398 10364
rect 7334 10304 7398 10308
rect 7414 10364 7478 10368
rect 7414 10308 7418 10364
rect 7418 10308 7474 10364
rect 7474 10308 7478 10364
rect 7414 10304 7478 10308
rect 7494 10364 7558 10368
rect 7494 10308 7498 10364
rect 7498 10308 7554 10364
rect 7554 10308 7558 10364
rect 7494 10304 7558 10308
rect 7574 10364 7638 10368
rect 7574 10308 7578 10364
rect 7578 10308 7634 10364
rect 7634 10308 7638 10364
rect 7574 10304 7638 10308
rect 9887 10364 9951 10368
rect 9887 10308 9891 10364
rect 9891 10308 9947 10364
rect 9947 10308 9951 10364
rect 9887 10304 9951 10308
rect 9967 10364 10031 10368
rect 9967 10308 9971 10364
rect 9971 10308 10027 10364
rect 10027 10308 10031 10364
rect 9967 10304 10031 10308
rect 10047 10364 10111 10368
rect 10047 10308 10051 10364
rect 10051 10308 10107 10364
rect 10107 10308 10111 10364
rect 10047 10304 10111 10308
rect 10127 10364 10191 10368
rect 10127 10308 10131 10364
rect 10131 10308 10187 10364
rect 10187 10308 10191 10364
rect 10127 10304 10191 10308
rect 3504 9820 3568 9824
rect 3504 9764 3508 9820
rect 3508 9764 3564 9820
rect 3564 9764 3568 9820
rect 3504 9760 3568 9764
rect 3584 9820 3648 9824
rect 3584 9764 3588 9820
rect 3588 9764 3644 9820
rect 3644 9764 3648 9820
rect 3584 9760 3648 9764
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 6057 9820 6121 9824
rect 6057 9764 6061 9820
rect 6061 9764 6117 9820
rect 6117 9764 6121 9820
rect 6057 9760 6121 9764
rect 6137 9820 6201 9824
rect 6137 9764 6141 9820
rect 6141 9764 6197 9820
rect 6197 9764 6201 9820
rect 6137 9760 6201 9764
rect 6217 9820 6281 9824
rect 6217 9764 6221 9820
rect 6221 9764 6277 9820
rect 6277 9764 6281 9820
rect 6217 9760 6281 9764
rect 6297 9820 6361 9824
rect 6297 9764 6301 9820
rect 6301 9764 6357 9820
rect 6357 9764 6361 9820
rect 6297 9760 6361 9764
rect 8610 9820 8674 9824
rect 8610 9764 8614 9820
rect 8614 9764 8670 9820
rect 8670 9764 8674 9820
rect 8610 9760 8674 9764
rect 8690 9820 8754 9824
rect 8690 9764 8694 9820
rect 8694 9764 8750 9820
rect 8750 9764 8754 9820
rect 8690 9760 8754 9764
rect 8770 9820 8834 9824
rect 8770 9764 8774 9820
rect 8774 9764 8830 9820
rect 8830 9764 8834 9820
rect 8770 9760 8834 9764
rect 8850 9820 8914 9824
rect 8850 9764 8854 9820
rect 8854 9764 8910 9820
rect 8910 9764 8914 9820
rect 8850 9760 8914 9764
rect 11163 9820 11227 9824
rect 11163 9764 11167 9820
rect 11167 9764 11223 9820
rect 11223 9764 11227 9820
rect 11163 9760 11227 9764
rect 11243 9820 11307 9824
rect 11243 9764 11247 9820
rect 11247 9764 11303 9820
rect 11303 9764 11307 9820
rect 11243 9760 11307 9764
rect 11323 9820 11387 9824
rect 11323 9764 11327 9820
rect 11327 9764 11383 9820
rect 11383 9764 11387 9820
rect 11323 9760 11387 9764
rect 11403 9820 11467 9824
rect 11403 9764 11407 9820
rect 11407 9764 11463 9820
rect 11463 9764 11467 9820
rect 11403 9760 11467 9764
rect 2228 9276 2292 9280
rect 2228 9220 2232 9276
rect 2232 9220 2288 9276
rect 2288 9220 2292 9276
rect 2228 9216 2292 9220
rect 2308 9276 2372 9280
rect 2308 9220 2312 9276
rect 2312 9220 2368 9276
rect 2368 9220 2372 9276
rect 2308 9216 2372 9220
rect 2388 9276 2452 9280
rect 2388 9220 2392 9276
rect 2392 9220 2448 9276
rect 2448 9220 2452 9276
rect 2388 9216 2452 9220
rect 2468 9276 2532 9280
rect 2468 9220 2472 9276
rect 2472 9220 2528 9276
rect 2528 9220 2532 9276
rect 2468 9216 2532 9220
rect 4781 9276 4845 9280
rect 4781 9220 4785 9276
rect 4785 9220 4841 9276
rect 4841 9220 4845 9276
rect 4781 9216 4845 9220
rect 4861 9276 4925 9280
rect 4861 9220 4865 9276
rect 4865 9220 4921 9276
rect 4921 9220 4925 9276
rect 4861 9216 4925 9220
rect 4941 9276 5005 9280
rect 4941 9220 4945 9276
rect 4945 9220 5001 9276
rect 5001 9220 5005 9276
rect 4941 9216 5005 9220
rect 5021 9276 5085 9280
rect 5021 9220 5025 9276
rect 5025 9220 5081 9276
rect 5081 9220 5085 9276
rect 5021 9216 5085 9220
rect 7334 9276 7398 9280
rect 7334 9220 7338 9276
rect 7338 9220 7394 9276
rect 7394 9220 7398 9276
rect 7334 9216 7398 9220
rect 7414 9276 7478 9280
rect 7414 9220 7418 9276
rect 7418 9220 7474 9276
rect 7474 9220 7478 9276
rect 7414 9216 7478 9220
rect 7494 9276 7558 9280
rect 7494 9220 7498 9276
rect 7498 9220 7554 9276
rect 7554 9220 7558 9276
rect 7494 9216 7558 9220
rect 7574 9276 7638 9280
rect 7574 9220 7578 9276
rect 7578 9220 7634 9276
rect 7634 9220 7638 9276
rect 7574 9216 7638 9220
rect 9887 9276 9951 9280
rect 9887 9220 9891 9276
rect 9891 9220 9947 9276
rect 9947 9220 9951 9276
rect 9887 9216 9951 9220
rect 9967 9276 10031 9280
rect 9967 9220 9971 9276
rect 9971 9220 10027 9276
rect 10027 9220 10031 9276
rect 9967 9216 10031 9220
rect 10047 9276 10111 9280
rect 10047 9220 10051 9276
rect 10051 9220 10107 9276
rect 10107 9220 10111 9276
rect 10047 9216 10111 9220
rect 10127 9276 10191 9280
rect 10127 9220 10131 9276
rect 10131 9220 10187 9276
rect 10187 9220 10191 9276
rect 10127 9216 10191 9220
rect 3504 8732 3568 8736
rect 3504 8676 3508 8732
rect 3508 8676 3564 8732
rect 3564 8676 3568 8732
rect 3504 8672 3568 8676
rect 3584 8732 3648 8736
rect 3584 8676 3588 8732
rect 3588 8676 3644 8732
rect 3644 8676 3648 8732
rect 3584 8672 3648 8676
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 6057 8732 6121 8736
rect 6057 8676 6061 8732
rect 6061 8676 6117 8732
rect 6117 8676 6121 8732
rect 6057 8672 6121 8676
rect 6137 8732 6201 8736
rect 6137 8676 6141 8732
rect 6141 8676 6197 8732
rect 6197 8676 6201 8732
rect 6137 8672 6201 8676
rect 6217 8732 6281 8736
rect 6217 8676 6221 8732
rect 6221 8676 6277 8732
rect 6277 8676 6281 8732
rect 6217 8672 6281 8676
rect 6297 8732 6361 8736
rect 6297 8676 6301 8732
rect 6301 8676 6357 8732
rect 6357 8676 6361 8732
rect 6297 8672 6361 8676
rect 8610 8732 8674 8736
rect 8610 8676 8614 8732
rect 8614 8676 8670 8732
rect 8670 8676 8674 8732
rect 8610 8672 8674 8676
rect 8690 8732 8754 8736
rect 8690 8676 8694 8732
rect 8694 8676 8750 8732
rect 8750 8676 8754 8732
rect 8690 8672 8754 8676
rect 8770 8732 8834 8736
rect 8770 8676 8774 8732
rect 8774 8676 8830 8732
rect 8830 8676 8834 8732
rect 8770 8672 8834 8676
rect 8850 8732 8914 8736
rect 8850 8676 8854 8732
rect 8854 8676 8910 8732
rect 8910 8676 8914 8732
rect 8850 8672 8914 8676
rect 11163 8732 11227 8736
rect 11163 8676 11167 8732
rect 11167 8676 11223 8732
rect 11223 8676 11227 8732
rect 11163 8672 11227 8676
rect 11243 8732 11307 8736
rect 11243 8676 11247 8732
rect 11247 8676 11303 8732
rect 11303 8676 11307 8732
rect 11243 8672 11307 8676
rect 11323 8732 11387 8736
rect 11323 8676 11327 8732
rect 11327 8676 11383 8732
rect 11383 8676 11387 8732
rect 11323 8672 11387 8676
rect 11403 8732 11467 8736
rect 11403 8676 11407 8732
rect 11407 8676 11463 8732
rect 11463 8676 11467 8732
rect 11403 8672 11467 8676
rect 2228 8188 2292 8192
rect 2228 8132 2232 8188
rect 2232 8132 2288 8188
rect 2288 8132 2292 8188
rect 2228 8128 2292 8132
rect 2308 8188 2372 8192
rect 2308 8132 2312 8188
rect 2312 8132 2368 8188
rect 2368 8132 2372 8188
rect 2308 8128 2372 8132
rect 2388 8188 2452 8192
rect 2388 8132 2392 8188
rect 2392 8132 2448 8188
rect 2448 8132 2452 8188
rect 2388 8128 2452 8132
rect 2468 8188 2532 8192
rect 2468 8132 2472 8188
rect 2472 8132 2528 8188
rect 2528 8132 2532 8188
rect 2468 8128 2532 8132
rect 4781 8188 4845 8192
rect 4781 8132 4785 8188
rect 4785 8132 4841 8188
rect 4841 8132 4845 8188
rect 4781 8128 4845 8132
rect 4861 8188 4925 8192
rect 4861 8132 4865 8188
rect 4865 8132 4921 8188
rect 4921 8132 4925 8188
rect 4861 8128 4925 8132
rect 4941 8188 5005 8192
rect 4941 8132 4945 8188
rect 4945 8132 5001 8188
rect 5001 8132 5005 8188
rect 4941 8128 5005 8132
rect 5021 8188 5085 8192
rect 5021 8132 5025 8188
rect 5025 8132 5081 8188
rect 5081 8132 5085 8188
rect 5021 8128 5085 8132
rect 7334 8188 7398 8192
rect 7334 8132 7338 8188
rect 7338 8132 7394 8188
rect 7394 8132 7398 8188
rect 7334 8128 7398 8132
rect 7414 8188 7478 8192
rect 7414 8132 7418 8188
rect 7418 8132 7474 8188
rect 7474 8132 7478 8188
rect 7414 8128 7478 8132
rect 7494 8188 7558 8192
rect 7494 8132 7498 8188
rect 7498 8132 7554 8188
rect 7554 8132 7558 8188
rect 7494 8128 7558 8132
rect 7574 8188 7638 8192
rect 7574 8132 7578 8188
rect 7578 8132 7634 8188
rect 7634 8132 7638 8188
rect 7574 8128 7638 8132
rect 9887 8188 9951 8192
rect 9887 8132 9891 8188
rect 9891 8132 9947 8188
rect 9947 8132 9951 8188
rect 9887 8128 9951 8132
rect 9967 8188 10031 8192
rect 9967 8132 9971 8188
rect 9971 8132 10027 8188
rect 10027 8132 10031 8188
rect 9967 8128 10031 8132
rect 10047 8188 10111 8192
rect 10047 8132 10051 8188
rect 10051 8132 10107 8188
rect 10107 8132 10111 8188
rect 10047 8128 10111 8132
rect 10127 8188 10191 8192
rect 10127 8132 10131 8188
rect 10131 8132 10187 8188
rect 10187 8132 10191 8188
rect 10127 8128 10191 8132
rect 3504 7644 3568 7648
rect 3504 7588 3508 7644
rect 3508 7588 3564 7644
rect 3564 7588 3568 7644
rect 3504 7584 3568 7588
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 6057 7644 6121 7648
rect 6057 7588 6061 7644
rect 6061 7588 6117 7644
rect 6117 7588 6121 7644
rect 6057 7584 6121 7588
rect 6137 7644 6201 7648
rect 6137 7588 6141 7644
rect 6141 7588 6197 7644
rect 6197 7588 6201 7644
rect 6137 7584 6201 7588
rect 6217 7644 6281 7648
rect 6217 7588 6221 7644
rect 6221 7588 6277 7644
rect 6277 7588 6281 7644
rect 6217 7584 6281 7588
rect 6297 7644 6361 7648
rect 6297 7588 6301 7644
rect 6301 7588 6357 7644
rect 6357 7588 6361 7644
rect 6297 7584 6361 7588
rect 8610 7644 8674 7648
rect 8610 7588 8614 7644
rect 8614 7588 8670 7644
rect 8670 7588 8674 7644
rect 8610 7584 8674 7588
rect 8690 7644 8754 7648
rect 8690 7588 8694 7644
rect 8694 7588 8750 7644
rect 8750 7588 8754 7644
rect 8690 7584 8754 7588
rect 8770 7644 8834 7648
rect 8770 7588 8774 7644
rect 8774 7588 8830 7644
rect 8830 7588 8834 7644
rect 8770 7584 8834 7588
rect 8850 7644 8914 7648
rect 8850 7588 8854 7644
rect 8854 7588 8910 7644
rect 8910 7588 8914 7644
rect 8850 7584 8914 7588
rect 11163 7644 11227 7648
rect 11163 7588 11167 7644
rect 11167 7588 11223 7644
rect 11223 7588 11227 7644
rect 11163 7584 11227 7588
rect 11243 7644 11307 7648
rect 11243 7588 11247 7644
rect 11247 7588 11303 7644
rect 11303 7588 11307 7644
rect 11243 7584 11307 7588
rect 11323 7644 11387 7648
rect 11323 7588 11327 7644
rect 11327 7588 11383 7644
rect 11383 7588 11387 7644
rect 11323 7584 11387 7588
rect 11403 7644 11467 7648
rect 11403 7588 11407 7644
rect 11407 7588 11463 7644
rect 11463 7588 11467 7644
rect 11403 7584 11467 7588
rect 2228 7100 2292 7104
rect 2228 7044 2232 7100
rect 2232 7044 2288 7100
rect 2288 7044 2292 7100
rect 2228 7040 2292 7044
rect 2308 7100 2372 7104
rect 2308 7044 2312 7100
rect 2312 7044 2368 7100
rect 2368 7044 2372 7100
rect 2308 7040 2372 7044
rect 2388 7100 2452 7104
rect 2388 7044 2392 7100
rect 2392 7044 2448 7100
rect 2448 7044 2452 7100
rect 2388 7040 2452 7044
rect 2468 7100 2532 7104
rect 2468 7044 2472 7100
rect 2472 7044 2528 7100
rect 2528 7044 2532 7100
rect 2468 7040 2532 7044
rect 4781 7100 4845 7104
rect 4781 7044 4785 7100
rect 4785 7044 4841 7100
rect 4841 7044 4845 7100
rect 4781 7040 4845 7044
rect 4861 7100 4925 7104
rect 4861 7044 4865 7100
rect 4865 7044 4921 7100
rect 4921 7044 4925 7100
rect 4861 7040 4925 7044
rect 4941 7100 5005 7104
rect 4941 7044 4945 7100
rect 4945 7044 5001 7100
rect 5001 7044 5005 7100
rect 4941 7040 5005 7044
rect 5021 7100 5085 7104
rect 5021 7044 5025 7100
rect 5025 7044 5081 7100
rect 5081 7044 5085 7100
rect 5021 7040 5085 7044
rect 7334 7100 7398 7104
rect 7334 7044 7338 7100
rect 7338 7044 7394 7100
rect 7394 7044 7398 7100
rect 7334 7040 7398 7044
rect 7414 7100 7478 7104
rect 7414 7044 7418 7100
rect 7418 7044 7474 7100
rect 7474 7044 7478 7100
rect 7414 7040 7478 7044
rect 7494 7100 7558 7104
rect 7494 7044 7498 7100
rect 7498 7044 7554 7100
rect 7554 7044 7558 7100
rect 7494 7040 7558 7044
rect 7574 7100 7638 7104
rect 7574 7044 7578 7100
rect 7578 7044 7634 7100
rect 7634 7044 7638 7100
rect 7574 7040 7638 7044
rect 9887 7100 9951 7104
rect 9887 7044 9891 7100
rect 9891 7044 9947 7100
rect 9947 7044 9951 7100
rect 9887 7040 9951 7044
rect 9967 7100 10031 7104
rect 9967 7044 9971 7100
rect 9971 7044 10027 7100
rect 10027 7044 10031 7100
rect 9967 7040 10031 7044
rect 10047 7100 10111 7104
rect 10047 7044 10051 7100
rect 10051 7044 10107 7100
rect 10107 7044 10111 7100
rect 10047 7040 10111 7044
rect 10127 7100 10191 7104
rect 10127 7044 10131 7100
rect 10131 7044 10187 7100
rect 10187 7044 10191 7100
rect 10127 7040 10191 7044
rect 3504 6556 3568 6560
rect 3504 6500 3508 6556
rect 3508 6500 3564 6556
rect 3564 6500 3568 6556
rect 3504 6496 3568 6500
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 6057 6556 6121 6560
rect 6057 6500 6061 6556
rect 6061 6500 6117 6556
rect 6117 6500 6121 6556
rect 6057 6496 6121 6500
rect 6137 6556 6201 6560
rect 6137 6500 6141 6556
rect 6141 6500 6197 6556
rect 6197 6500 6201 6556
rect 6137 6496 6201 6500
rect 6217 6556 6281 6560
rect 6217 6500 6221 6556
rect 6221 6500 6277 6556
rect 6277 6500 6281 6556
rect 6217 6496 6281 6500
rect 6297 6556 6361 6560
rect 6297 6500 6301 6556
rect 6301 6500 6357 6556
rect 6357 6500 6361 6556
rect 6297 6496 6361 6500
rect 8610 6556 8674 6560
rect 8610 6500 8614 6556
rect 8614 6500 8670 6556
rect 8670 6500 8674 6556
rect 8610 6496 8674 6500
rect 8690 6556 8754 6560
rect 8690 6500 8694 6556
rect 8694 6500 8750 6556
rect 8750 6500 8754 6556
rect 8690 6496 8754 6500
rect 8770 6556 8834 6560
rect 8770 6500 8774 6556
rect 8774 6500 8830 6556
rect 8830 6500 8834 6556
rect 8770 6496 8834 6500
rect 8850 6556 8914 6560
rect 8850 6500 8854 6556
rect 8854 6500 8910 6556
rect 8910 6500 8914 6556
rect 8850 6496 8914 6500
rect 11163 6556 11227 6560
rect 11163 6500 11167 6556
rect 11167 6500 11223 6556
rect 11223 6500 11227 6556
rect 11163 6496 11227 6500
rect 11243 6556 11307 6560
rect 11243 6500 11247 6556
rect 11247 6500 11303 6556
rect 11303 6500 11307 6556
rect 11243 6496 11307 6500
rect 11323 6556 11387 6560
rect 11323 6500 11327 6556
rect 11327 6500 11383 6556
rect 11383 6500 11387 6556
rect 11323 6496 11387 6500
rect 11403 6556 11467 6560
rect 11403 6500 11407 6556
rect 11407 6500 11463 6556
rect 11463 6500 11467 6556
rect 11403 6496 11467 6500
rect 2228 6012 2292 6016
rect 2228 5956 2232 6012
rect 2232 5956 2288 6012
rect 2288 5956 2292 6012
rect 2228 5952 2292 5956
rect 2308 6012 2372 6016
rect 2308 5956 2312 6012
rect 2312 5956 2368 6012
rect 2368 5956 2372 6012
rect 2308 5952 2372 5956
rect 2388 6012 2452 6016
rect 2388 5956 2392 6012
rect 2392 5956 2448 6012
rect 2448 5956 2452 6012
rect 2388 5952 2452 5956
rect 2468 6012 2532 6016
rect 2468 5956 2472 6012
rect 2472 5956 2528 6012
rect 2528 5956 2532 6012
rect 2468 5952 2532 5956
rect 4781 6012 4845 6016
rect 4781 5956 4785 6012
rect 4785 5956 4841 6012
rect 4841 5956 4845 6012
rect 4781 5952 4845 5956
rect 4861 6012 4925 6016
rect 4861 5956 4865 6012
rect 4865 5956 4921 6012
rect 4921 5956 4925 6012
rect 4861 5952 4925 5956
rect 4941 6012 5005 6016
rect 4941 5956 4945 6012
rect 4945 5956 5001 6012
rect 5001 5956 5005 6012
rect 4941 5952 5005 5956
rect 5021 6012 5085 6016
rect 5021 5956 5025 6012
rect 5025 5956 5081 6012
rect 5081 5956 5085 6012
rect 5021 5952 5085 5956
rect 7334 6012 7398 6016
rect 7334 5956 7338 6012
rect 7338 5956 7394 6012
rect 7394 5956 7398 6012
rect 7334 5952 7398 5956
rect 7414 6012 7478 6016
rect 7414 5956 7418 6012
rect 7418 5956 7474 6012
rect 7474 5956 7478 6012
rect 7414 5952 7478 5956
rect 7494 6012 7558 6016
rect 7494 5956 7498 6012
rect 7498 5956 7554 6012
rect 7554 5956 7558 6012
rect 7494 5952 7558 5956
rect 7574 6012 7638 6016
rect 7574 5956 7578 6012
rect 7578 5956 7634 6012
rect 7634 5956 7638 6012
rect 7574 5952 7638 5956
rect 9887 6012 9951 6016
rect 9887 5956 9891 6012
rect 9891 5956 9947 6012
rect 9947 5956 9951 6012
rect 9887 5952 9951 5956
rect 9967 6012 10031 6016
rect 9967 5956 9971 6012
rect 9971 5956 10027 6012
rect 10027 5956 10031 6012
rect 9967 5952 10031 5956
rect 10047 6012 10111 6016
rect 10047 5956 10051 6012
rect 10051 5956 10107 6012
rect 10107 5956 10111 6012
rect 10047 5952 10111 5956
rect 10127 6012 10191 6016
rect 10127 5956 10131 6012
rect 10131 5956 10187 6012
rect 10187 5956 10191 6012
rect 10127 5952 10191 5956
rect 3504 5468 3568 5472
rect 3504 5412 3508 5468
rect 3508 5412 3564 5468
rect 3564 5412 3568 5468
rect 3504 5408 3568 5412
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 6057 5468 6121 5472
rect 6057 5412 6061 5468
rect 6061 5412 6117 5468
rect 6117 5412 6121 5468
rect 6057 5408 6121 5412
rect 6137 5468 6201 5472
rect 6137 5412 6141 5468
rect 6141 5412 6197 5468
rect 6197 5412 6201 5468
rect 6137 5408 6201 5412
rect 6217 5468 6281 5472
rect 6217 5412 6221 5468
rect 6221 5412 6277 5468
rect 6277 5412 6281 5468
rect 6217 5408 6281 5412
rect 6297 5468 6361 5472
rect 6297 5412 6301 5468
rect 6301 5412 6357 5468
rect 6357 5412 6361 5468
rect 6297 5408 6361 5412
rect 8610 5468 8674 5472
rect 8610 5412 8614 5468
rect 8614 5412 8670 5468
rect 8670 5412 8674 5468
rect 8610 5408 8674 5412
rect 8690 5468 8754 5472
rect 8690 5412 8694 5468
rect 8694 5412 8750 5468
rect 8750 5412 8754 5468
rect 8690 5408 8754 5412
rect 8770 5468 8834 5472
rect 8770 5412 8774 5468
rect 8774 5412 8830 5468
rect 8830 5412 8834 5468
rect 8770 5408 8834 5412
rect 8850 5468 8914 5472
rect 8850 5412 8854 5468
rect 8854 5412 8910 5468
rect 8910 5412 8914 5468
rect 8850 5408 8914 5412
rect 11163 5468 11227 5472
rect 11163 5412 11167 5468
rect 11167 5412 11223 5468
rect 11223 5412 11227 5468
rect 11163 5408 11227 5412
rect 11243 5468 11307 5472
rect 11243 5412 11247 5468
rect 11247 5412 11303 5468
rect 11303 5412 11307 5468
rect 11243 5408 11307 5412
rect 11323 5468 11387 5472
rect 11323 5412 11327 5468
rect 11327 5412 11383 5468
rect 11383 5412 11387 5468
rect 11323 5408 11387 5412
rect 11403 5468 11467 5472
rect 11403 5412 11407 5468
rect 11407 5412 11463 5468
rect 11463 5412 11467 5468
rect 11403 5408 11467 5412
rect 2228 4924 2292 4928
rect 2228 4868 2232 4924
rect 2232 4868 2288 4924
rect 2288 4868 2292 4924
rect 2228 4864 2292 4868
rect 2308 4924 2372 4928
rect 2308 4868 2312 4924
rect 2312 4868 2368 4924
rect 2368 4868 2372 4924
rect 2308 4864 2372 4868
rect 2388 4924 2452 4928
rect 2388 4868 2392 4924
rect 2392 4868 2448 4924
rect 2448 4868 2452 4924
rect 2388 4864 2452 4868
rect 2468 4924 2532 4928
rect 2468 4868 2472 4924
rect 2472 4868 2528 4924
rect 2528 4868 2532 4924
rect 2468 4864 2532 4868
rect 4781 4924 4845 4928
rect 4781 4868 4785 4924
rect 4785 4868 4841 4924
rect 4841 4868 4845 4924
rect 4781 4864 4845 4868
rect 4861 4924 4925 4928
rect 4861 4868 4865 4924
rect 4865 4868 4921 4924
rect 4921 4868 4925 4924
rect 4861 4864 4925 4868
rect 4941 4924 5005 4928
rect 4941 4868 4945 4924
rect 4945 4868 5001 4924
rect 5001 4868 5005 4924
rect 4941 4864 5005 4868
rect 5021 4924 5085 4928
rect 5021 4868 5025 4924
rect 5025 4868 5081 4924
rect 5081 4868 5085 4924
rect 5021 4864 5085 4868
rect 7334 4924 7398 4928
rect 7334 4868 7338 4924
rect 7338 4868 7394 4924
rect 7394 4868 7398 4924
rect 7334 4864 7398 4868
rect 7414 4924 7478 4928
rect 7414 4868 7418 4924
rect 7418 4868 7474 4924
rect 7474 4868 7478 4924
rect 7414 4864 7478 4868
rect 7494 4924 7558 4928
rect 7494 4868 7498 4924
rect 7498 4868 7554 4924
rect 7554 4868 7558 4924
rect 7494 4864 7558 4868
rect 7574 4924 7638 4928
rect 7574 4868 7578 4924
rect 7578 4868 7634 4924
rect 7634 4868 7638 4924
rect 7574 4864 7638 4868
rect 9887 4924 9951 4928
rect 9887 4868 9891 4924
rect 9891 4868 9947 4924
rect 9947 4868 9951 4924
rect 9887 4864 9951 4868
rect 9967 4924 10031 4928
rect 9967 4868 9971 4924
rect 9971 4868 10027 4924
rect 10027 4868 10031 4924
rect 9967 4864 10031 4868
rect 10047 4924 10111 4928
rect 10047 4868 10051 4924
rect 10051 4868 10107 4924
rect 10107 4868 10111 4924
rect 10047 4864 10111 4868
rect 10127 4924 10191 4928
rect 10127 4868 10131 4924
rect 10131 4868 10187 4924
rect 10187 4868 10191 4924
rect 10127 4864 10191 4868
rect 3504 4380 3568 4384
rect 3504 4324 3508 4380
rect 3508 4324 3564 4380
rect 3564 4324 3568 4380
rect 3504 4320 3568 4324
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 6057 4380 6121 4384
rect 6057 4324 6061 4380
rect 6061 4324 6117 4380
rect 6117 4324 6121 4380
rect 6057 4320 6121 4324
rect 6137 4380 6201 4384
rect 6137 4324 6141 4380
rect 6141 4324 6197 4380
rect 6197 4324 6201 4380
rect 6137 4320 6201 4324
rect 6217 4380 6281 4384
rect 6217 4324 6221 4380
rect 6221 4324 6277 4380
rect 6277 4324 6281 4380
rect 6217 4320 6281 4324
rect 6297 4380 6361 4384
rect 6297 4324 6301 4380
rect 6301 4324 6357 4380
rect 6357 4324 6361 4380
rect 6297 4320 6361 4324
rect 8610 4380 8674 4384
rect 8610 4324 8614 4380
rect 8614 4324 8670 4380
rect 8670 4324 8674 4380
rect 8610 4320 8674 4324
rect 8690 4380 8754 4384
rect 8690 4324 8694 4380
rect 8694 4324 8750 4380
rect 8750 4324 8754 4380
rect 8690 4320 8754 4324
rect 8770 4380 8834 4384
rect 8770 4324 8774 4380
rect 8774 4324 8830 4380
rect 8830 4324 8834 4380
rect 8770 4320 8834 4324
rect 8850 4380 8914 4384
rect 8850 4324 8854 4380
rect 8854 4324 8910 4380
rect 8910 4324 8914 4380
rect 8850 4320 8914 4324
rect 11163 4380 11227 4384
rect 11163 4324 11167 4380
rect 11167 4324 11223 4380
rect 11223 4324 11227 4380
rect 11163 4320 11227 4324
rect 11243 4380 11307 4384
rect 11243 4324 11247 4380
rect 11247 4324 11303 4380
rect 11303 4324 11307 4380
rect 11243 4320 11307 4324
rect 11323 4380 11387 4384
rect 11323 4324 11327 4380
rect 11327 4324 11383 4380
rect 11383 4324 11387 4380
rect 11323 4320 11387 4324
rect 11403 4380 11467 4384
rect 11403 4324 11407 4380
rect 11407 4324 11463 4380
rect 11463 4324 11467 4380
rect 11403 4320 11467 4324
rect 2228 3836 2292 3840
rect 2228 3780 2232 3836
rect 2232 3780 2288 3836
rect 2288 3780 2292 3836
rect 2228 3776 2292 3780
rect 2308 3836 2372 3840
rect 2308 3780 2312 3836
rect 2312 3780 2368 3836
rect 2368 3780 2372 3836
rect 2308 3776 2372 3780
rect 2388 3836 2452 3840
rect 2388 3780 2392 3836
rect 2392 3780 2448 3836
rect 2448 3780 2452 3836
rect 2388 3776 2452 3780
rect 2468 3836 2532 3840
rect 2468 3780 2472 3836
rect 2472 3780 2528 3836
rect 2528 3780 2532 3836
rect 2468 3776 2532 3780
rect 4781 3836 4845 3840
rect 4781 3780 4785 3836
rect 4785 3780 4841 3836
rect 4841 3780 4845 3836
rect 4781 3776 4845 3780
rect 4861 3836 4925 3840
rect 4861 3780 4865 3836
rect 4865 3780 4921 3836
rect 4921 3780 4925 3836
rect 4861 3776 4925 3780
rect 4941 3836 5005 3840
rect 4941 3780 4945 3836
rect 4945 3780 5001 3836
rect 5001 3780 5005 3836
rect 4941 3776 5005 3780
rect 5021 3836 5085 3840
rect 5021 3780 5025 3836
rect 5025 3780 5081 3836
rect 5081 3780 5085 3836
rect 5021 3776 5085 3780
rect 7334 3836 7398 3840
rect 7334 3780 7338 3836
rect 7338 3780 7394 3836
rect 7394 3780 7398 3836
rect 7334 3776 7398 3780
rect 7414 3836 7478 3840
rect 7414 3780 7418 3836
rect 7418 3780 7474 3836
rect 7474 3780 7478 3836
rect 7414 3776 7478 3780
rect 7494 3836 7558 3840
rect 7494 3780 7498 3836
rect 7498 3780 7554 3836
rect 7554 3780 7558 3836
rect 7494 3776 7558 3780
rect 7574 3836 7638 3840
rect 7574 3780 7578 3836
rect 7578 3780 7634 3836
rect 7634 3780 7638 3836
rect 7574 3776 7638 3780
rect 9887 3836 9951 3840
rect 9887 3780 9891 3836
rect 9891 3780 9947 3836
rect 9947 3780 9951 3836
rect 9887 3776 9951 3780
rect 9967 3836 10031 3840
rect 9967 3780 9971 3836
rect 9971 3780 10027 3836
rect 10027 3780 10031 3836
rect 9967 3776 10031 3780
rect 10047 3836 10111 3840
rect 10047 3780 10051 3836
rect 10051 3780 10107 3836
rect 10107 3780 10111 3836
rect 10047 3776 10111 3780
rect 10127 3836 10191 3840
rect 10127 3780 10131 3836
rect 10131 3780 10187 3836
rect 10187 3780 10191 3836
rect 10127 3776 10191 3780
rect 3504 3292 3568 3296
rect 3504 3236 3508 3292
rect 3508 3236 3564 3292
rect 3564 3236 3568 3292
rect 3504 3232 3568 3236
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 6057 3292 6121 3296
rect 6057 3236 6061 3292
rect 6061 3236 6117 3292
rect 6117 3236 6121 3292
rect 6057 3232 6121 3236
rect 6137 3292 6201 3296
rect 6137 3236 6141 3292
rect 6141 3236 6197 3292
rect 6197 3236 6201 3292
rect 6137 3232 6201 3236
rect 6217 3292 6281 3296
rect 6217 3236 6221 3292
rect 6221 3236 6277 3292
rect 6277 3236 6281 3292
rect 6217 3232 6281 3236
rect 6297 3292 6361 3296
rect 6297 3236 6301 3292
rect 6301 3236 6357 3292
rect 6357 3236 6361 3292
rect 6297 3232 6361 3236
rect 8610 3292 8674 3296
rect 8610 3236 8614 3292
rect 8614 3236 8670 3292
rect 8670 3236 8674 3292
rect 8610 3232 8674 3236
rect 8690 3292 8754 3296
rect 8690 3236 8694 3292
rect 8694 3236 8750 3292
rect 8750 3236 8754 3292
rect 8690 3232 8754 3236
rect 8770 3292 8834 3296
rect 8770 3236 8774 3292
rect 8774 3236 8830 3292
rect 8830 3236 8834 3292
rect 8770 3232 8834 3236
rect 8850 3292 8914 3296
rect 8850 3236 8854 3292
rect 8854 3236 8910 3292
rect 8910 3236 8914 3292
rect 8850 3232 8914 3236
rect 11163 3292 11227 3296
rect 11163 3236 11167 3292
rect 11167 3236 11223 3292
rect 11223 3236 11227 3292
rect 11163 3232 11227 3236
rect 11243 3292 11307 3296
rect 11243 3236 11247 3292
rect 11247 3236 11303 3292
rect 11303 3236 11307 3292
rect 11243 3232 11307 3236
rect 11323 3292 11387 3296
rect 11323 3236 11327 3292
rect 11327 3236 11383 3292
rect 11383 3236 11387 3292
rect 11323 3232 11387 3236
rect 11403 3292 11467 3296
rect 11403 3236 11407 3292
rect 11407 3236 11463 3292
rect 11463 3236 11467 3292
rect 11403 3232 11467 3236
rect 2228 2748 2292 2752
rect 2228 2692 2232 2748
rect 2232 2692 2288 2748
rect 2288 2692 2292 2748
rect 2228 2688 2292 2692
rect 2308 2748 2372 2752
rect 2308 2692 2312 2748
rect 2312 2692 2368 2748
rect 2368 2692 2372 2748
rect 2308 2688 2372 2692
rect 2388 2748 2452 2752
rect 2388 2692 2392 2748
rect 2392 2692 2448 2748
rect 2448 2692 2452 2748
rect 2388 2688 2452 2692
rect 2468 2748 2532 2752
rect 2468 2692 2472 2748
rect 2472 2692 2528 2748
rect 2528 2692 2532 2748
rect 2468 2688 2532 2692
rect 4781 2748 4845 2752
rect 4781 2692 4785 2748
rect 4785 2692 4841 2748
rect 4841 2692 4845 2748
rect 4781 2688 4845 2692
rect 4861 2748 4925 2752
rect 4861 2692 4865 2748
rect 4865 2692 4921 2748
rect 4921 2692 4925 2748
rect 4861 2688 4925 2692
rect 4941 2748 5005 2752
rect 4941 2692 4945 2748
rect 4945 2692 5001 2748
rect 5001 2692 5005 2748
rect 4941 2688 5005 2692
rect 5021 2748 5085 2752
rect 5021 2692 5025 2748
rect 5025 2692 5081 2748
rect 5081 2692 5085 2748
rect 5021 2688 5085 2692
rect 7334 2748 7398 2752
rect 7334 2692 7338 2748
rect 7338 2692 7394 2748
rect 7394 2692 7398 2748
rect 7334 2688 7398 2692
rect 7414 2748 7478 2752
rect 7414 2692 7418 2748
rect 7418 2692 7474 2748
rect 7474 2692 7478 2748
rect 7414 2688 7478 2692
rect 7494 2748 7558 2752
rect 7494 2692 7498 2748
rect 7498 2692 7554 2748
rect 7554 2692 7558 2748
rect 7494 2688 7558 2692
rect 7574 2748 7638 2752
rect 7574 2692 7578 2748
rect 7578 2692 7634 2748
rect 7634 2692 7638 2748
rect 7574 2688 7638 2692
rect 9887 2748 9951 2752
rect 9887 2692 9891 2748
rect 9891 2692 9947 2748
rect 9947 2692 9951 2748
rect 9887 2688 9951 2692
rect 9967 2748 10031 2752
rect 9967 2692 9971 2748
rect 9971 2692 10027 2748
rect 10027 2692 10031 2748
rect 9967 2688 10031 2692
rect 10047 2748 10111 2752
rect 10047 2692 10051 2748
rect 10051 2692 10107 2748
rect 10107 2692 10111 2748
rect 10047 2688 10111 2692
rect 10127 2748 10191 2752
rect 10127 2692 10131 2748
rect 10131 2692 10187 2748
rect 10187 2692 10191 2748
rect 10127 2688 10191 2692
rect 3504 2204 3568 2208
rect 3504 2148 3508 2204
rect 3508 2148 3564 2204
rect 3564 2148 3568 2204
rect 3504 2144 3568 2148
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 6057 2204 6121 2208
rect 6057 2148 6061 2204
rect 6061 2148 6117 2204
rect 6117 2148 6121 2204
rect 6057 2144 6121 2148
rect 6137 2204 6201 2208
rect 6137 2148 6141 2204
rect 6141 2148 6197 2204
rect 6197 2148 6201 2204
rect 6137 2144 6201 2148
rect 6217 2204 6281 2208
rect 6217 2148 6221 2204
rect 6221 2148 6277 2204
rect 6277 2148 6281 2204
rect 6217 2144 6281 2148
rect 6297 2204 6361 2208
rect 6297 2148 6301 2204
rect 6301 2148 6357 2204
rect 6357 2148 6361 2204
rect 6297 2144 6361 2148
rect 8610 2204 8674 2208
rect 8610 2148 8614 2204
rect 8614 2148 8670 2204
rect 8670 2148 8674 2204
rect 8610 2144 8674 2148
rect 8690 2204 8754 2208
rect 8690 2148 8694 2204
rect 8694 2148 8750 2204
rect 8750 2148 8754 2204
rect 8690 2144 8754 2148
rect 8770 2204 8834 2208
rect 8770 2148 8774 2204
rect 8774 2148 8830 2204
rect 8830 2148 8834 2204
rect 8770 2144 8834 2148
rect 8850 2204 8914 2208
rect 8850 2148 8854 2204
rect 8854 2148 8910 2204
rect 8910 2148 8914 2204
rect 8850 2144 8914 2148
rect 11163 2204 11227 2208
rect 11163 2148 11167 2204
rect 11167 2148 11223 2204
rect 11223 2148 11227 2204
rect 11163 2144 11227 2148
rect 11243 2204 11307 2208
rect 11243 2148 11247 2204
rect 11247 2148 11303 2204
rect 11303 2148 11307 2204
rect 11243 2144 11307 2148
rect 11323 2204 11387 2208
rect 11323 2148 11327 2204
rect 11327 2148 11383 2204
rect 11383 2148 11387 2204
rect 11323 2144 11387 2148
rect 11403 2204 11467 2208
rect 11403 2148 11407 2204
rect 11407 2148 11463 2204
rect 11463 2148 11467 2204
rect 11403 2144 11467 2148
<< metal4 >>
rect 3496 12086 3816 12128
rect 2220 11456 2540 12016
rect 2220 11392 2228 11456
rect 2292 11392 2308 11456
rect 2372 11392 2388 11456
rect 2452 11392 2468 11456
rect 2532 11392 2540 11456
rect 2220 10862 2540 11392
rect 2220 10626 2262 10862
rect 2498 10626 2540 10862
rect 2220 10368 2540 10626
rect 2220 10304 2228 10368
rect 2292 10304 2308 10368
rect 2372 10304 2388 10368
rect 2452 10304 2468 10368
rect 2532 10304 2540 10368
rect 2220 9280 2540 10304
rect 2220 9216 2228 9280
rect 2292 9216 2308 9280
rect 2372 9216 2388 9280
rect 2452 9216 2468 9280
rect 2532 9216 2540 9280
rect 2220 8414 2540 9216
rect 2220 8192 2262 8414
rect 2498 8192 2540 8414
rect 2220 8128 2228 8192
rect 2292 8128 2308 8178
rect 2372 8128 2388 8178
rect 2452 8128 2468 8178
rect 2532 8128 2540 8192
rect 2220 7104 2540 8128
rect 2220 7040 2228 7104
rect 2292 7040 2308 7104
rect 2372 7040 2388 7104
rect 2452 7040 2468 7104
rect 2532 7040 2540 7104
rect 2220 6016 2540 7040
rect 2220 5952 2228 6016
rect 2292 5966 2308 6016
rect 2372 5966 2388 6016
rect 2452 5966 2468 6016
rect 2532 5952 2540 6016
rect 2220 5730 2262 5952
rect 2498 5730 2540 5952
rect 2220 4928 2540 5730
rect 2220 4864 2228 4928
rect 2292 4864 2308 4928
rect 2372 4864 2388 4928
rect 2452 4864 2468 4928
rect 2532 4864 2540 4928
rect 2220 3840 2540 4864
rect 2220 3776 2228 3840
rect 2292 3776 2308 3840
rect 2372 3776 2388 3840
rect 2452 3776 2468 3840
rect 2532 3776 2540 3840
rect 2220 3518 2540 3776
rect 2220 3282 2262 3518
rect 2498 3282 2540 3518
rect 2220 2752 2540 3282
rect 2220 2688 2228 2752
rect 2292 2688 2308 2752
rect 2372 2688 2388 2752
rect 2452 2688 2468 2752
rect 2532 2688 2540 2752
rect 2220 2128 2540 2688
rect 3496 12000 3538 12086
rect 3774 12000 3816 12086
rect 6049 12086 6369 12128
rect 3496 11936 3504 12000
rect 3808 11936 3816 12000
rect 3496 11850 3538 11936
rect 3774 11850 3816 11936
rect 3496 10912 3816 11850
rect 3496 10848 3504 10912
rect 3568 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3816 10912
rect 3496 9824 3816 10848
rect 3496 9760 3504 9824
rect 3568 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3816 9824
rect 3496 9638 3816 9760
rect 3496 9402 3538 9638
rect 3774 9402 3816 9638
rect 3496 8736 3816 9402
rect 3496 8672 3504 8736
rect 3568 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3816 8736
rect 3496 7648 3816 8672
rect 3496 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3816 7648
rect 3496 7190 3816 7584
rect 3496 6954 3538 7190
rect 3774 6954 3816 7190
rect 3496 6560 3816 6954
rect 3496 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3816 6560
rect 3496 5472 3816 6496
rect 3496 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3816 5472
rect 3496 4742 3816 5408
rect 3496 4506 3538 4742
rect 3774 4506 3816 4742
rect 3496 4384 3816 4506
rect 3496 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3816 4384
rect 3496 3296 3816 4320
rect 3496 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3816 3296
rect 3496 2208 3816 3232
rect 3496 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3816 2208
rect 3496 2128 3816 2144
rect 4773 11456 5093 12016
rect 4773 11392 4781 11456
rect 4845 11392 4861 11456
rect 4925 11392 4941 11456
rect 5005 11392 5021 11456
rect 5085 11392 5093 11456
rect 4773 10862 5093 11392
rect 4773 10626 4815 10862
rect 5051 10626 5093 10862
rect 4773 10368 5093 10626
rect 4773 10304 4781 10368
rect 4845 10304 4861 10368
rect 4925 10304 4941 10368
rect 5005 10304 5021 10368
rect 5085 10304 5093 10368
rect 4773 9280 5093 10304
rect 4773 9216 4781 9280
rect 4845 9216 4861 9280
rect 4925 9216 4941 9280
rect 5005 9216 5021 9280
rect 5085 9216 5093 9280
rect 4773 8414 5093 9216
rect 4773 8192 4815 8414
rect 5051 8192 5093 8414
rect 4773 8128 4781 8192
rect 4845 8128 4861 8178
rect 4925 8128 4941 8178
rect 5005 8128 5021 8178
rect 5085 8128 5093 8192
rect 4773 7104 5093 8128
rect 4773 7040 4781 7104
rect 4845 7040 4861 7104
rect 4925 7040 4941 7104
rect 5005 7040 5021 7104
rect 5085 7040 5093 7104
rect 4773 6016 5093 7040
rect 4773 5952 4781 6016
rect 4845 5966 4861 6016
rect 4925 5966 4941 6016
rect 5005 5966 5021 6016
rect 5085 5952 5093 6016
rect 4773 5730 4815 5952
rect 5051 5730 5093 5952
rect 4773 4928 5093 5730
rect 4773 4864 4781 4928
rect 4845 4864 4861 4928
rect 4925 4864 4941 4928
rect 5005 4864 5021 4928
rect 5085 4864 5093 4928
rect 4773 3840 5093 4864
rect 4773 3776 4781 3840
rect 4845 3776 4861 3840
rect 4925 3776 4941 3840
rect 5005 3776 5021 3840
rect 5085 3776 5093 3840
rect 4773 3518 5093 3776
rect 4773 3282 4815 3518
rect 5051 3282 5093 3518
rect 4773 2752 5093 3282
rect 4773 2688 4781 2752
rect 4845 2688 4861 2752
rect 4925 2688 4941 2752
rect 5005 2688 5021 2752
rect 5085 2688 5093 2752
rect 4773 2128 5093 2688
rect 6049 12000 6091 12086
rect 6327 12000 6369 12086
rect 8602 12086 8922 12128
rect 6049 11936 6057 12000
rect 6361 11936 6369 12000
rect 6049 11850 6091 11936
rect 6327 11850 6369 11936
rect 6049 10912 6369 11850
rect 6049 10848 6057 10912
rect 6121 10848 6137 10912
rect 6201 10848 6217 10912
rect 6281 10848 6297 10912
rect 6361 10848 6369 10912
rect 6049 9824 6369 10848
rect 6049 9760 6057 9824
rect 6121 9760 6137 9824
rect 6201 9760 6217 9824
rect 6281 9760 6297 9824
rect 6361 9760 6369 9824
rect 6049 9638 6369 9760
rect 6049 9402 6091 9638
rect 6327 9402 6369 9638
rect 6049 8736 6369 9402
rect 6049 8672 6057 8736
rect 6121 8672 6137 8736
rect 6201 8672 6217 8736
rect 6281 8672 6297 8736
rect 6361 8672 6369 8736
rect 6049 7648 6369 8672
rect 6049 7584 6057 7648
rect 6121 7584 6137 7648
rect 6201 7584 6217 7648
rect 6281 7584 6297 7648
rect 6361 7584 6369 7648
rect 6049 7190 6369 7584
rect 6049 6954 6091 7190
rect 6327 6954 6369 7190
rect 6049 6560 6369 6954
rect 6049 6496 6057 6560
rect 6121 6496 6137 6560
rect 6201 6496 6217 6560
rect 6281 6496 6297 6560
rect 6361 6496 6369 6560
rect 6049 5472 6369 6496
rect 6049 5408 6057 5472
rect 6121 5408 6137 5472
rect 6201 5408 6217 5472
rect 6281 5408 6297 5472
rect 6361 5408 6369 5472
rect 6049 4742 6369 5408
rect 6049 4506 6091 4742
rect 6327 4506 6369 4742
rect 6049 4384 6369 4506
rect 6049 4320 6057 4384
rect 6121 4320 6137 4384
rect 6201 4320 6217 4384
rect 6281 4320 6297 4384
rect 6361 4320 6369 4384
rect 6049 3296 6369 4320
rect 6049 3232 6057 3296
rect 6121 3232 6137 3296
rect 6201 3232 6217 3296
rect 6281 3232 6297 3296
rect 6361 3232 6369 3296
rect 6049 2208 6369 3232
rect 6049 2144 6057 2208
rect 6121 2144 6137 2208
rect 6201 2144 6217 2208
rect 6281 2144 6297 2208
rect 6361 2144 6369 2208
rect 6049 2128 6369 2144
rect 7326 11456 7646 12016
rect 7326 11392 7334 11456
rect 7398 11392 7414 11456
rect 7478 11392 7494 11456
rect 7558 11392 7574 11456
rect 7638 11392 7646 11456
rect 7326 10862 7646 11392
rect 7326 10626 7368 10862
rect 7604 10626 7646 10862
rect 7326 10368 7646 10626
rect 7326 10304 7334 10368
rect 7398 10304 7414 10368
rect 7478 10304 7494 10368
rect 7558 10304 7574 10368
rect 7638 10304 7646 10368
rect 7326 9280 7646 10304
rect 7326 9216 7334 9280
rect 7398 9216 7414 9280
rect 7478 9216 7494 9280
rect 7558 9216 7574 9280
rect 7638 9216 7646 9280
rect 7326 8414 7646 9216
rect 7326 8192 7368 8414
rect 7604 8192 7646 8414
rect 7326 8128 7334 8192
rect 7398 8128 7414 8178
rect 7478 8128 7494 8178
rect 7558 8128 7574 8178
rect 7638 8128 7646 8192
rect 7326 7104 7646 8128
rect 7326 7040 7334 7104
rect 7398 7040 7414 7104
rect 7478 7040 7494 7104
rect 7558 7040 7574 7104
rect 7638 7040 7646 7104
rect 7326 6016 7646 7040
rect 7326 5952 7334 6016
rect 7398 5966 7414 6016
rect 7478 5966 7494 6016
rect 7558 5966 7574 6016
rect 7638 5952 7646 6016
rect 7326 5730 7368 5952
rect 7604 5730 7646 5952
rect 7326 4928 7646 5730
rect 7326 4864 7334 4928
rect 7398 4864 7414 4928
rect 7478 4864 7494 4928
rect 7558 4864 7574 4928
rect 7638 4864 7646 4928
rect 7326 3840 7646 4864
rect 7326 3776 7334 3840
rect 7398 3776 7414 3840
rect 7478 3776 7494 3840
rect 7558 3776 7574 3840
rect 7638 3776 7646 3840
rect 7326 3518 7646 3776
rect 7326 3282 7368 3518
rect 7604 3282 7646 3518
rect 7326 2752 7646 3282
rect 7326 2688 7334 2752
rect 7398 2688 7414 2752
rect 7478 2688 7494 2752
rect 7558 2688 7574 2752
rect 7638 2688 7646 2752
rect 7326 2128 7646 2688
rect 8602 12000 8644 12086
rect 8880 12000 8922 12086
rect 11155 12086 11475 12128
rect 8602 11936 8610 12000
rect 8914 11936 8922 12000
rect 8602 11850 8644 11936
rect 8880 11850 8922 11936
rect 8602 10912 8922 11850
rect 8602 10848 8610 10912
rect 8674 10848 8690 10912
rect 8754 10848 8770 10912
rect 8834 10848 8850 10912
rect 8914 10848 8922 10912
rect 8602 9824 8922 10848
rect 8602 9760 8610 9824
rect 8674 9760 8690 9824
rect 8754 9760 8770 9824
rect 8834 9760 8850 9824
rect 8914 9760 8922 9824
rect 8602 9638 8922 9760
rect 8602 9402 8644 9638
rect 8880 9402 8922 9638
rect 8602 8736 8922 9402
rect 8602 8672 8610 8736
rect 8674 8672 8690 8736
rect 8754 8672 8770 8736
rect 8834 8672 8850 8736
rect 8914 8672 8922 8736
rect 8602 7648 8922 8672
rect 8602 7584 8610 7648
rect 8674 7584 8690 7648
rect 8754 7584 8770 7648
rect 8834 7584 8850 7648
rect 8914 7584 8922 7648
rect 8602 7190 8922 7584
rect 8602 6954 8644 7190
rect 8880 6954 8922 7190
rect 8602 6560 8922 6954
rect 8602 6496 8610 6560
rect 8674 6496 8690 6560
rect 8754 6496 8770 6560
rect 8834 6496 8850 6560
rect 8914 6496 8922 6560
rect 8602 5472 8922 6496
rect 8602 5408 8610 5472
rect 8674 5408 8690 5472
rect 8754 5408 8770 5472
rect 8834 5408 8850 5472
rect 8914 5408 8922 5472
rect 8602 4742 8922 5408
rect 8602 4506 8644 4742
rect 8880 4506 8922 4742
rect 8602 4384 8922 4506
rect 8602 4320 8610 4384
rect 8674 4320 8690 4384
rect 8754 4320 8770 4384
rect 8834 4320 8850 4384
rect 8914 4320 8922 4384
rect 8602 3296 8922 4320
rect 8602 3232 8610 3296
rect 8674 3232 8690 3296
rect 8754 3232 8770 3296
rect 8834 3232 8850 3296
rect 8914 3232 8922 3296
rect 8602 2208 8922 3232
rect 8602 2144 8610 2208
rect 8674 2144 8690 2208
rect 8754 2144 8770 2208
rect 8834 2144 8850 2208
rect 8914 2144 8922 2208
rect 8602 2128 8922 2144
rect 9879 11456 10199 12016
rect 9879 11392 9887 11456
rect 9951 11392 9967 11456
rect 10031 11392 10047 11456
rect 10111 11392 10127 11456
rect 10191 11392 10199 11456
rect 9879 10862 10199 11392
rect 9879 10626 9921 10862
rect 10157 10626 10199 10862
rect 9879 10368 10199 10626
rect 9879 10304 9887 10368
rect 9951 10304 9967 10368
rect 10031 10304 10047 10368
rect 10111 10304 10127 10368
rect 10191 10304 10199 10368
rect 9879 9280 10199 10304
rect 9879 9216 9887 9280
rect 9951 9216 9967 9280
rect 10031 9216 10047 9280
rect 10111 9216 10127 9280
rect 10191 9216 10199 9280
rect 9879 8414 10199 9216
rect 9879 8192 9921 8414
rect 10157 8192 10199 8414
rect 9879 8128 9887 8192
rect 9951 8128 9967 8178
rect 10031 8128 10047 8178
rect 10111 8128 10127 8178
rect 10191 8128 10199 8192
rect 9879 7104 10199 8128
rect 9879 7040 9887 7104
rect 9951 7040 9967 7104
rect 10031 7040 10047 7104
rect 10111 7040 10127 7104
rect 10191 7040 10199 7104
rect 9879 6016 10199 7040
rect 9879 5952 9887 6016
rect 9951 5966 9967 6016
rect 10031 5966 10047 6016
rect 10111 5966 10127 6016
rect 10191 5952 10199 6016
rect 9879 5730 9921 5952
rect 10157 5730 10199 5952
rect 9879 4928 10199 5730
rect 9879 4864 9887 4928
rect 9951 4864 9967 4928
rect 10031 4864 10047 4928
rect 10111 4864 10127 4928
rect 10191 4864 10199 4928
rect 9879 3840 10199 4864
rect 9879 3776 9887 3840
rect 9951 3776 9967 3840
rect 10031 3776 10047 3840
rect 10111 3776 10127 3840
rect 10191 3776 10199 3840
rect 9879 3518 10199 3776
rect 9879 3282 9921 3518
rect 10157 3282 10199 3518
rect 9879 2752 10199 3282
rect 9879 2688 9887 2752
rect 9951 2688 9967 2752
rect 10031 2688 10047 2752
rect 10111 2688 10127 2752
rect 10191 2688 10199 2752
rect 9879 2128 10199 2688
rect 11155 12000 11197 12086
rect 11433 12000 11475 12086
rect 11155 11936 11163 12000
rect 11467 11936 11475 12000
rect 11155 11850 11197 11936
rect 11433 11850 11475 11936
rect 11155 10912 11475 11850
rect 11155 10848 11163 10912
rect 11227 10848 11243 10912
rect 11307 10848 11323 10912
rect 11387 10848 11403 10912
rect 11467 10848 11475 10912
rect 11155 9824 11475 10848
rect 11155 9760 11163 9824
rect 11227 9760 11243 9824
rect 11307 9760 11323 9824
rect 11387 9760 11403 9824
rect 11467 9760 11475 9824
rect 11155 9638 11475 9760
rect 11155 9402 11197 9638
rect 11433 9402 11475 9638
rect 11155 8736 11475 9402
rect 11155 8672 11163 8736
rect 11227 8672 11243 8736
rect 11307 8672 11323 8736
rect 11387 8672 11403 8736
rect 11467 8672 11475 8736
rect 11155 7648 11475 8672
rect 11155 7584 11163 7648
rect 11227 7584 11243 7648
rect 11307 7584 11323 7648
rect 11387 7584 11403 7648
rect 11467 7584 11475 7648
rect 11155 7190 11475 7584
rect 11155 6954 11197 7190
rect 11433 6954 11475 7190
rect 11155 6560 11475 6954
rect 11155 6496 11163 6560
rect 11227 6496 11243 6560
rect 11307 6496 11323 6560
rect 11387 6496 11403 6560
rect 11467 6496 11475 6560
rect 11155 5472 11475 6496
rect 11155 5408 11163 5472
rect 11227 5408 11243 5472
rect 11307 5408 11323 5472
rect 11387 5408 11403 5472
rect 11467 5408 11475 5472
rect 11155 4742 11475 5408
rect 11155 4506 11197 4742
rect 11433 4506 11475 4742
rect 11155 4384 11475 4506
rect 11155 4320 11163 4384
rect 11227 4320 11243 4384
rect 11307 4320 11323 4384
rect 11387 4320 11403 4384
rect 11467 4320 11475 4384
rect 11155 3296 11475 4320
rect 11155 3232 11163 3296
rect 11227 3232 11243 3296
rect 11307 3232 11323 3296
rect 11387 3232 11403 3296
rect 11467 3232 11475 3296
rect 11155 2208 11475 3232
rect 11155 2144 11163 2208
rect 11227 2144 11243 2208
rect 11307 2144 11323 2208
rect 11387 2144 11403 2208
rect 11467 2144 11475 2208
rect 11155 2128 11475 2144
<< via4 >>
rect 2262 10626 2498 10862
rect 2262 8192 2498 8414
rect 2262 8178 2292 8192
rect 2292 8178 2308 8192
rect 2308 8178 2372 8192
rect 2372 8178 2388 8192
rect 2388 8178 2452 8192
rect 2452 8178 2468 8192
rect 2468 8178 2498 8192
rect 2262 5952 2292 5966
rect 2292 5952 2308 5966
rect 2308 5952 2372 5966
rect 2372 5952 2388 5966
rect 2388 5952 2452 5966
rect 2452 5952 2468 5966
rect 2468 5952 2498 5966
rect 2262 5730 2498 5952
rect 2262 3282 2498 3518
rect 3538 12000 3774 12086
rect 3538 11936 3568 12000
rect 3568 11936 3584 12000
rect 3584 11936 3648 12000
rect 3648 11936 3664 12000
rect 3664 11936 3728 12000
rect 3728 11936 3744 12000
rect 3744 11936 3774 12000
rect 3538 11850 3774 11936
rect 3538 9402 3774 9638
rect 3538 6954 3774 7190
rect 3538 4506 3774 4742
rect 4815 10626 5051 10862
rect 4815 8192 5051 8414
rect 4815 8178 4845 8192
rect 4845 8178 4861 8192
rect 4861 8178 4925 8192
rect 4925 8178 4941 8192
rect 4941 8178 5005 8192
rect 5005 8178 5021 8192
rect 5021 8178 5051 8192
rect 4815 5952 4845 5966
rect 4845 5952 4861 5966
rect 4861 5952 4925 5966
rect 4925 5952 4941 5966
rect 4941 5952 5005 5966
rect 5005 5952 5021 5966
rect 5021 5952 5051 5966
rect 4815 5730 5051 5952
rect 4815 3282 5051 3518
rect 6091 12000 6327 12086
rect 6091 11936 6121 12000
rect 6121 11936 6137 12000
rect 6137 11936 6201 12000
rect 6201 11936 6217 12000
rect 6217 11936 6281 12000
rect 6281 11936 6297 12000
rect 6297 11936 6327 12000
rect 6091 11850 6327 11936
rect 6091 9402 6327 9638
rect 6091 6954 6327 7190
rect 6091 4506 6327 4742
rect 7368 10626 7604 10862
rect 7368 8192 7604 8414
rect 7368 8178 7398 8192
rect 7398 8178 7414 8192
rect 7414 8178 7478 8192
rect 7478 8178 7494 8192
rect 7494 8178 7558 8192
rect 7558 8178 7574 8192
rect 7574 8178 7604 8192
rect 7368 5952 7398 5966
rect 7398 5952 7414 5966
rect 7414 5952 7478 5966
rect 7478 5952 7494 5966
rect 7494 5952 7558 5966
rect 7558 5952 7574 5966
rect 7574 5952 7604 5966
rect 7368 5730 7604 5952
rect 7368 3282 7604 3518
rect 8644 12000 8880 12086
rect 8644 11936 8674 12000
rect 8674 11936 8690 12000
rect 8690 11936 8754 12000
rect 8754 11936 8770 12000
rect 8770 11936 8834 12000
rect 8834 11936 8850 12000
rect 8850 11936 8880 12000
rect 8644 11850 8880 11936
rect 8644 9402 8880 9638
rect 8644 6954 8880 7190
rect 8644 4506 8880 4742
rect 9921 10626 10157 10862
rect 9921 8192 10157 8414
rect 9921 8178 9951 8192
rect 9951 8178 9967 8192
rect 9967 8178 10031 8192
rect 10031 8178 10047 8192
rect 10047 8178 10111 8192
rect 10111 8178 10127 8192
rect 10127 8178 10157 8192
rect 9921 5952 9951 5966
rect 9951 5952 9967 5966
rect 9967 5952 10031 5966
rect 10031 5952 10047 5966
rect 10047 5952 10111 5966
rect 10111 5952 10127 5966
rect 10127 5952 10157 5966
rect 9921 5730 10157 5952
rect 9921 3282 10157 3518
rect 11197 12000 11433 12086
rect 11197 11936 11227 12000
rect 11227 11936 11243 12000
rect 11243 11936 11307 12000
rect 11307 11936 11323 12000
rect 11323 11936 11387 12000
rect 11387 11936 11403 12000
rect 11403 11936 11433 12000
rect 11197 11850 11433 11936
rect 11197 9402 11433 9638
rect 11197 6954 11433 7190
rect 11197 4506 11433 4742
<< metal5 >>
rect 1056 12086 11475 12128
rect 1056 11850 3538 12086
rect 3774 11850 6091 12086
rect 6327 11850 8644 12086
rect 8880 11850 11197 12086
rect 11433 11850 11475 12086
rect 1056 11808 11475 11850
rect 1056 10862 11364 10904
rect 1056 10626 2262 10862
rect 2498 10626 4815 10862
rect 5051 10626 7368 10862
rect 7604 10626 9921 10862
rect 10157 10626 11364 10862
rect 1056 10584 11364 10626
rect 1056 9638 11475 9680
rect 1056 9402 3538 9638
rect 3774 9402 6091 9638
rect 6327 9402 8644 9638
rect 8880 9402 11197 9638
rect 11433 9402 11475 9638
rect 1056 9360 11475 9402
rect 1056 8414 11364 8456
rect 1056 8178 2262 8414
rect 2498 8178 4815 8414
rect 5051 8178 7368 8414
rect 7604 8178 9921 8414
rect 10157 8178 11364 8414
rect 1056 8136 11364 8178
rect 1056 7190 11475 7232
rect 1056 6954 3538 7190
rect 3774 6954 6091 7190
rect 6327 6954 8644 7190
rect 8880 6954 11197 7190
rect 11433 6954 11475 7190
rect 1056 6912 11475 6954
rect 1056 5966 11364 6008
rect 1056 5730 2262 5966
rect 2498 5730 4815 5966
rect 5051 5730 7368 5966
rect 7604 5730 9921 5966
rect 10157 5730 11364 5966
rect 1056 5688 11364 5730
rect 1056 4742 11475 4784
rect 1056 4506 3538 4742
rect 3774 4506 6091 4742
rect 6327 4506 8644 4742
rect 8880 4506 11197 4742
rect 11433 4506 11475 4742
rect 1056 4464 11475 4506
rect 1056 3518 11364 3560
rect 1056 3282 2262 3518
rect 2498 3282 4815 3518
rect 5051 3282 7368 3518
rect 7604 3282 9921 3518
rect 10157 3282 11364 3518
rect 1056 3240 11364 3282
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1660669191
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1660669191
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1660669191
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1660669191
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1660669191
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1660669191
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1660669191
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1660669191
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1660669191
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1660669191
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1660669191
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1660669191
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1660669191
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1660669191
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1660669191
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1660669191
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1660669191
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp 1660669191
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1660669191
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1660669191
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1660669191
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1660669191
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1660669191
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_56
timestamp 1660669191
transform 1 0 6256 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_68
timestamp 1660669191
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1660669191
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1660669191
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1660669191
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1660669191
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_105
timestamp 1660669191
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1660669191
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1660669191
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1660669191
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1660669191
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1660669191
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1660669191
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1660669191
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1660669191
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_76
timestamp 1660669191
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_88
timestamp 1660669191
transform 1 0 9200 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_100
timestamp 1660669191
transform 1 0 10304 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1660669191
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1660669191
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1660669191
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1660669191
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1660669191
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1660669191
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1660669191
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1660669191
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1660669191
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1660669191
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp 1660669191
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_105
timestamp 1660669191
transform 1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1660669191
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1660669191
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1660669191
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1660669191
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1660669191
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1660669191
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1660669191
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1660669191
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1660669191
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1660669191
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp 1660669191
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1660669191
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1660669191
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1660669191
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1660669191
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1660669191
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1660669191
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1660669191
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1660669191
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1660669191
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1660669191
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1660669191
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1660669191
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1660669191
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1660669191
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1660669191
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1660669191
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1660669191
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1660669191
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1660669191
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1660669191
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1660669191
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1660669191
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp 1660669191
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1660669191
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1660669191
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1660669191
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1660669191
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1660669191
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1660669191
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1660669191
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1660669191
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1660669191
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1660669191
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1660669191
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_105
timestamp 1660669191
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1660669191
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1660669191
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1660669191
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1660669191
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1660669191
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1660669191
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1660669191
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1660669191
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1660669191
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1660669191
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp 1660669191
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1660669191
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1660669191
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1660669191
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1660669191
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1660669191
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1660669191
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1660669191
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1660669191
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1660669191
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1660669191
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_101
timestamp 1660669191
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_107
timestamp 1660669191
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1660669191
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1660669191
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1660669191
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1660669191
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1660669191
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1660669191
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1660669191
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_62
timestamp 1660669191
transform 1 0 6808 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_74
timestamp 1660669191
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_82
timestamp 1660669191
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_105
timestamp 1660669191
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1660669191
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1660669191
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1660669191
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1660669191
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1660669191
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1660669191
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_51
timestamp 1660669191
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_63
timestamp 1660669191
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1660669191
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1660669191
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1660669191
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1660669191
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_105
timestamp 1660669191
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1660669191
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1660669191
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1660669191
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_30
timestamp 1660669191
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1660669191
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1660669191
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1660669191
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1660669191
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1660669191
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_94
timestamp 1660669191
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1660669191
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1660669191
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1660669191
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1660669191
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1660669191
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1660669191
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1660669191
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1660669191
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1660669191
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1660669191
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1660669191
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1660669191
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1660669191
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1660669191
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1660669191
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1660669191
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1660669191
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1660669191
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1660669191
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1660669191
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1660669191
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_105
timestamp 1660669191
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1660669191
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1660669191
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1660669191
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1660669191
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1660669191
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1660669191
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1660669191
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1660669191
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1660669191
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1660669191
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1660669191
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_105
timestamp 1660669191
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1660669191
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1660669191
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_21
timestamp 1660669191
transform 1 0 3036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1660669191
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1660669191
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1660669191
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1660669191
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1660669191
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1660669191
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1660669191
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_81
timestamp 1660669191
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_85
timestamp 1660669191
transform 1 0 8924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1660669191
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1660669191
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1660669191
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1660669191
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1660669191
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1660669191
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1660669191
transform -1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1660669191
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1660669191
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1660669191
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1660669191
transform -1 0 11316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1660669191
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1660669191
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1660669191
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1660669191
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1660669191
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1660669191
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1660669191
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1660669191
transform -1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1660669191
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1660669191
transform -1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1660669191
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1660669191
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1660669191
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1660669191
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1660669191
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1660669191
transform -1 0 11316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1660669191
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1660669191
transform -1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1660669191
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1660669191
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1660669191
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1660669191
transform -1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1660669191
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1660669191
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1660669191
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1660669191
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1660669191
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1660669191
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1660669191
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1660669191
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1660669191
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1660669191
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1660669191
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1660669191
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1660669191
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1660669191
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1660669191
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1660669191
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1660669191
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1660669191
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1660669191
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1660669191
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1660669191
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1660669191
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1660669191
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1660669191
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1660669191
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1660669191
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1660669191
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1660669191
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1660669191
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1660669191
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1660669191
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1660669191
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1660669191
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1660669191
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1660669191
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 3128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _07_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 5520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 2484 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1660669191
transform -1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 1660669191
transform 1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1660669191
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1660669191
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1660669191
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 5244 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 10764 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform -1 0 9752 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1660669191
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1660669191
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1660669191
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1660669191
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1660669191
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1660669191
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1660669191
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1660669191
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1660669191
transform -1 0 4324 0 -1 11968
box -38 -48 406 592
<< labels >>
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 C
port 0 nsew signal input
flabel metal4 s 3496 2128 3816 12128 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 6049 2128 6369 12128 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8602 2128 8922 12128 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 11155 2128 11475 12128 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 4464 11475 4784 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 6912 11475 7232 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 9360 11475 9680 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 11808 11475 12128 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2220 2128 2540 12016 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 4773 2128 5093 12016 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 7326 2128 7646 12016 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 9879 2128 10199 12016 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 3240 11364 3560 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 5688 11364 6008 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 8136 11364 8456 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 10584 11364 10904 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 clk
port 3 nsew signal input
flabel metal2 s 9678 13852 9734 14652 0 FreeSans 224 90 0 0 light_farm[0]
port 4 nsew signal tristate
flabel metal3 s 11708 11568 12508 11688 0 FreeSans 480 0 0 0 light_farm[1]
port 5 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 light_farm[2]
port 6 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 light_highway[0]
port 7 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 light_highway[1]
port 8 nsew signal tristate
flabel metal2 s 3238 13852 3294 14652 0 FreeSans 224 90 0 0 light_highway[2]
port 9 nsew signal tristate
flabel metal3 s 11708 5448 12508 5568 0 FreeSans 480 0 0 0 rst_n
port 10 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12508 14652
<< end >>
